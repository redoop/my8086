module MyCPU8086(
  input         clock,
  input         reset,
  output [19:0] io_memAddr, // @[src/main/scala/cpu8086/CPU8086.scala 22:14]
  output [15:0] io_memDataOut, // @[src/main/scala/cpu8086/CPU8086.scala 22:14]
  input  [15:0] io_memDataIn, // @[src/main/scala/cpu8086/CPU8086.scala 22:14]
  output        io_memWrite, // @[src/main/scala/cpu8086/CPU8086.scala 22:14]
  output        io_memRead, // @[src/main/scala/cpu8086/CPU8086.scala 22:14]
  output        io_halt, // @[src/main/scala/cpu8086/CPU8086.scala 22:14]
  output [15:0] io_ax, // @[src/main/scala/cpu8086/CPU8086.scala 22:14]
  output [15:0] io_bx, // @[src/main/scala/cpu8086/CPU8086.scala 22:14]
  output [15:0] io_cx, // @[src/main/scala/cpu8086/CPU8086.scala 22:14]
  output [15:0] io_dx, // @[src/main/scala/cpu8086/CPU8086.scala 22:14]
  output [15:0] io_sp, // @[src/main/scala/cpu8086/CPU8086.scala 22:14]
  output [15:0] io_ip, // @[src/main/scala/cpu8086/CPU8086.scala 22:14]
  output [15:0] io_flags // @[src/main/scala/cpu8086/CPU8086.scala 22:14]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
`endif // RANDOMIZE_REG_INIT
  reg [15:0] ax; // @[src/main/scala/cpu8086/CPU8086.scala 40:19]
  reg [15:0] bx; // @[src/main/scala/cpu8086/CPU8086.scala 41:19]
  reg [15:0] cx; // @[src/main/scala/cpu8086/CPU8086.scala 42:19]
  reg [15:0] dx; // @[src/main/scala/cpu8086/CPU8086.scala 43:19]
  reg [15:0] sp; // @[src/main/scala/cpu8086/CPU8086.scala 44:19]
  reg [15:0] bp; // @[src/main/scala/cpu8086/CPU8086.scala 45:19]
  reg [15:0] si; // @[src/main/scala/cpu8086/CPU8086.scala 46:19]
  reg [15:0] di; // @[src/main/scala/cpu8086/CPU8086.scala 47:19]
  reg [15:0] ip; // @[src/main/scala/cpu8086/CPU8086.scala 56:19]
  reg [15:0] flags; // @[src/main/scala/cpu8086/CPU8086.scala 57:22]
  reg [2:0] state; // @[src/main/scala/cpu8086/CPU8086.scala 61:22]
  reg [15:0] instruction; // @[src/main/scala/cpu8086/CPU8086.scala 63:28]
  reg [15:0] memData; // @[src/main/scala/cpu8086/CPU8086.scala 64:24]
  wire [19:0] _GEN_787 = {{4'd0}, ip}; // @[src/main/scala/cpu8086/CPU8086.scala 139:27]
  wire [19:0] _io_memAddr_T_2 = 20'hffff0 + _GEN_787; // @[src/main/scala/cpu8086/CPU8086.scala 139:27]
  wire [15:0] _ip_T_1 = ip + 16'h2; // @[src/main/scala/cpu8086/CPU8086.scala 157:16]
  wire [7:0] opcode = instruction[15:8]; // @[src/main/scala/cpu8086/CPU8086.scala 162:31]
  wire [7:0] operand = instruction[7:0]; // @[src/main/scala/cpu8086/CPU8086.scala 163:32]
  wire [2:0] srcReg = operand[2:0]; // @[src/main/scala/cpu8086/CPU8086.scala 164:27]
  wire [2:0] dstReg = operand[5:3]; // @[src/main/scala/cpu8086/CPU8086.scala 165:27]
  wire  _srcVal_T = 3'h1 == srcReg; // @[src/main/scala/cpu8086/CPU8086.scala 97:27]
  wire [15:0] _srcVal_T_1 = 3'h1 == srcReg ? cx : ax; // @[src/main/scala/cpu8086/CPU8086.scala 97:27]
  wire  _srcVal_T_2 = 3'h2 == srcReg; // @[src/main/scala/cpu8086/CPU8086.scala 97:27]
  wire [15:0] _srcVal_T_3 = 3'h2 == srcReg ? dx : _srcVal_T_1; // @[src/main/scala/cpu8086/CPU8086.scala 97:27]
  wire  _srcVal_T_4 = 3'h3 == srcReg; // @[src/main/scala/cpu8086/CPU8086.scala 97:27]
  wire [15:0] _srcVal_T_5 = 3'h3 == srcReg ? bx : _srcVal_T_3; // @[src/main/scala/cpu8086/CPU8086.scala 97:27]
  wire  _srcVal_T_6 = 3'h4 == srcReg; // @[src/main/scala/cpu8086/CPU8086.scala 97:27]
  wire [15:0] _srcVal_T_7 = 3'h4 == srcReg ? sp : _srcVal_T_5; // @[src/main/scala/cpu8086/CPU8086.scala 97:27]
  wire  _srcVal_T_8 = 3'h5 == srcReg; // @[src/main/scala/cpu8086/CPU8086.scala 97:27]
  wire [15:0] _srcVal_T_9 = 3'h5 == srcReg ? bp : _srcVal_T_7; // @[src/main/scala/cpu8086/CPU8086.scala 97:27]
  wire  _srcVal_T_10 = 3'h6 == srcReg; // @[src/main/scala/cpu8086/CPU8086.scala 97:27]
  wire [15:0] _srcVal_T_11 = 3'h6 == srcReg ? si : _srcVal_T_9; // @[src/main/scala/cpu8086/CPU8086.scala 97:27]
  wire  _srcVal_T_12 = 3'h7 == srcReg; // @[src/main/scala/cpu8086/CPU8086.scala 97:27]
  wire [15:0] srcVal = 3'h7 == srcReg ? di : _srcVal_T_11; // @[src/main/scala/cpu8086/CPU8086.scala 97:27]
  wire  _T_4 = 3'h1 == dstReg; // @[src/main/scala/cpu8086/CPU8086.scala 110:21]
  wire  _T_5 = 3'h2 == dstReg; // @[src/main/scala/cpu8086/CPU8086.scala 110:21]
  wire  _T_6 = 3'h3 == dstReg; // @[src/main/scala/cpu8086/CPU8086.scala 110:21]
  wire  _T_7 = 3'h4 == dstReg; // @[src/main/scala/cpu8086/CPU8086.scala 110:21]
  wire  _T_8 = 3'h5 == dstReg; // @[src/main/scala/cpu8086/CPU8086.scala 110:21]
  wire  _T_9 = 3'h6 == dstReg; // @[src/main/scala/cpu8086/CPU8086.scala 110:21]
  wire  _T_10 = 3'h7 == dstReg; // @[src/main/scala/cpu8086/CPU8086.scala 110:21]
  wire [15:0] _GEN_0 = 3'h7 == dstReg ? srcVal : di; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 118:20 47:19]
  wire [15:0] _GEN_1 = 3'h6 == dstReg ? srcVal : si; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 117:20 46:19]
  wire [15:0] _GEN_2 = 3'h6 == dstReg ? di : _GEN_0; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 47:19]
  wire [15:0] _GEN_3 = 3'h5 == dstReg ? srcVal : bp; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 116:20 45:19]
  wire [15:0] _GEN_4 = 3'h5 == dstReg ? si : _GEN_1; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 46:19]
  wire [15:0] _GEN_5 = 3'h5 == dstReg ? di : _GEN_2; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 47:19]
  wire [15:0] _GEN_6 = 3'h4 == dstReg ? srcVal : sp; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 115:20 44:19]
  wire [15:0] _GEN_7 = 3'h4 == dstReg ? bp : _GEN_3; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 45:19]
  wire [15:0] _GEN_8 = 3'h4 == dstReg ? si : _GEN_4; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 46:19]
  wire [15:0] _GEN_9 = 3'h4 == dstReg ? di : _GEN_5; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 47:19]
  wire [15:0] _GEN_10 = 3'h3 == dstReg ? srcVal : bx; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 114:20 41:19]
  wire [15:0] _GEN_11 = 3'h3 == dstReg ? sp : _GEN_6; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 44:19]
  wire [15:0] _GEN_12 = 3'h3 == dstReg ? bp : _GEN_7; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 45:19]
  wire [15:0] _GEN_13 = 3'h3 == dstReg ? si : _GEN_8; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 46:19]
  wire [15:0] _GEN_14 = 3'h3 == dstReg ? di : _GEN_9; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 47:19]
  wire [15:0] _GEN_15 = 3'h2 == dstReg ? srcVal : dx; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 113:20 43:19]
  wire [15:0] _GEN_16 = 3'h2 == dstReg ? bx : _GEN_10; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 41:19]
  wire [15:0] _GEN_17 = 3'h2 == dstReg ? sp : _GEN_11; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 44:19]
  wire [15:0] _GEN_18 = 3'h2 == dstReg ? bp : _GEN_12; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 45:19]
  wire [15:0] _GEN_19 = 3'h2 == dstReg ? si : _GEN_13; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 46:19]
  wire [15:0] _GEN_20 = 3'h2 == dstReg ? di : _GEN_14; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 47:19]
  wire [15:0] _GEN_21 = 3'h1 == dstReg ? srcVal : cx; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 112:20 42:19]
  wire [15:0] _GEN_22 = 3'h1 == dstReg ? dx : _GEN_15; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 43:19]
  wire [15:0] _GEN_23 = 3'h1 == dstReg ? bx : _GEN_16; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 41:19]
  wire [15:0] _GEN_24 = 3'h1 == dstReg ? sp : _GEN_17; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 44:19]
  wire [15:0] _GEN_25 = 3'h1 == dstReg ? bp : _GEN_18; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 45:19]
  wire [15:0] _GEN_26 = 3'h1 == dstReg ? si : _GEN_19; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 46:19]
  wire [15:0] _GEN_27 = 3'h1 == dstReg ? di : _GEN_20; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 47:19]
  wire [15:0] _GEN_28 = 3'h0 == dstReg ? srcVal : ax; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 111:20 40:19]
  wire [15:0] _GEN_29 = 3'h0 == dstReg ? cx : _GEN_21; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 42:19]
  wire [15:0] _GEN_30 = 3'h0 == dstReg ? dx : _GEN_22; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 43:19]
  wire [15:0] _GEN_31 = 3'h0 == dstReg ? bx : _GEN_23; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 41:19]
  wire [15:0] _GEN_32 = 3'h0 == dstReg ? sp : _GEN_24; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 44:19]
  wire [15:0] _GEN_33 = 3'h0 == dstReg ? bp : _GEN_25; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 45:19]
  wire [15:0] _GEN_34 = 3'h0 == dstReg ? si : _GEN_26; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 46:19]
  wire [15:0] _GEN_35 = 3'h0 == dstReg ? di : _GEN_27; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 47:19]
  wire [15:0] _ax_T = {operand,8'h0}; // @[src/main/scala/cpu8086/CPU8086.scala 179:25]
  wire [15:0] _dst_T_1 = _T_4 ? cx : ax; // @[src/main/scala/cpu8086/CPU8086.scala 97:27]
  wire [15:0] _dst_T_3 = _T_5 ? dx : _dst_T_1; // @[src/main/scala/cpu8086/CPU8086.scala 97:27]
  wire [15:0] _dst_T_5 = _T_6 ? bx : _dst_T_3; // @[src/main/scala/cpu8086/CPU8086.scala 97:27]
  wire [15:0] _dst_T_7 = _T_7 ? sp : _dst_T_5; // @[src/main/scala/cpu8086/CPU8086.scala 97:27]
  wire [15:0] _dst_T_9 = _T_8 ? bp : _dst_T_7; // @[src/main/scala/cpu8086/CPU8086.scala 97:27]
  wire [15:0] _dst_T_11 = _T_9 ? si : _dst_T_9; // @[src/main/scala/cpu8086/CPU8086.scala 97:27]
  wire [15:0] dst = _T_10 ? di : _dst_T_11; // @[src/main/scala/cpu8086/CPU8086.scala 97:27]
  wire [16:0] result = dst + srcVal; // @[src/main/scala/cpu8086/CPU8086.scala 207:28]
  wire  carryOut = result[16]; // @[src/main/scala/cpu8086/CPU8086.scala 208:32]
  wire  overflow = dst[15] == srcVal[15] & dst[15] != result[15]; // @[src/main/scala/cpu8086/CPU8086.scala 209:48]
  wire [15:0] _GEN_36 = 3'h7 == dstReg ? result[15:0] : di; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 118:20 47:19]
  wire [15:0] _GEN_37 = 3'h6 == dstReg ? result[15:0] : si; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 117:20 46:19]
  wire [15:0] _GEN_38 = 3'h6 == dstReg ? di : _GEN_36; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 47:19]
  wire [15:0] _GEN_39 = 3'h5 == dstReg ? result[15:0] : bp; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 116:20 45:19]
  wire [15:0] _GEN_40 = 3'h5 == dstReg ? si : _GEN_37; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 46:19]
  wire [15:0] _GEN_41 = 3'h5 == dstReg ? di : _GEN_38; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 47:19]
  wire [15:0] _GEN_42 = 3'h4 == dstReg ? result[15:0] : sp; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 115:20 44:19]
  wire [15:0] _GEN_43 = 3'h4 == dstReg ? bp : _GEN_39; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 45:19]
  wire [15:0] _GEN_44 = 3'h4 == dstReg ? si : _GEN_40; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 46:19]
  wire [15:0] _GEN_45 = 3'h4 == dstReg ? di : _GEN_41; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 47:19]
  wire [15:0] _GEN_46 = 3'h3 == dstReg ? result[15:0] : bx; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 114:20 41:19]
  wire [15:0] _GEN_47 = 3'h3 == dstReg ? sp : _GEN_42; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 44:19]
  wire [15:0] _GEN_48 = 3'h3 == dstReg ? bp : _GEN_43; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 45:19]
  wire [15:0] _GEN_49 = 3'h3 == dstReg ? si : _GEN_44; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 46:19]
  wire [15:0] _GEN_50 = 3'h3 == dstReg ? di : _GEN_45; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 47:19]
  wire [15:0] _GEN_51 = 3'h2 == dstReg ? result[15:0] : dx; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 113:20 43:19]
  wire [15:0] _GEN_52 = 3'h2 == dstReg ? bx : _GEN_46; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 41:19]
  wire [15:0] _GEN_53 = 3'h2 == dstReg ? sp : _GEN_47; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 44:19]
  wire [15:0] _GEN_54 = 3'h2 == dstReg ? bp : _GEN_48; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 45:19]
  wire [15:0] _GEN_55 = 3'h2 == dstReg ? si : _GEN_49; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 46:19]
  wire [15:0] _GEN_56 = 3'h2 == dstReg ? di : _GEN_50; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 47:19]
  wire [15:0] _GEN_57 = 3'h1 == dstReg ? result[15:0] : cx; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 112:20 42:19]
  wire [15:0] _GEN_58 = 3'h1 == dstReg ? dx : _GEN_51; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 43:19]
  wire [15:0] _GEN_59 = 3'h1 == dstReg ? bx : _GEN_52; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 41:19]
  wire [15:0] _GEN_60 = 3'h1 == dstReg ? sp : _GEN_53; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 44:19]
  wire [15:0] _GEN_61 = 3'h1 == dstReg ? bp : _GEN_54; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 45:19]
  wire [15:0] _GEN_62 = 3'h1 == dstReg ? si : _GEN_55; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 46:19]
  wire [15:0] _GEN_63 = 3'h1 == dstReg ? di : _GEN_56; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 47:19]
  wire [15:0] _GEN_64 = 3'h0 == dstReg ? result[15:0] : ax; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 111:20 40:19]
  wire [15:0] _GEN_65 = 3'h0 == dstReg ? cx : _GEN_57; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 42:19]
  wire [15:0] _GEN_66 = 3'h0 == dstReg ? dx : _GEN_58; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 43:19]
  wire [15:0] _GEN_67 = 3'h0 == dstReg ? bx : _GEN_59; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 41:19]
  wire [15:0] _GEN_68 = 3'h0 == dstReg ? sp : _GEN_60; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 44:19]
  wire [15:0] _GEN_69 = 3'h0 == dstReg ? bp : _GEN_61; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 45:19]
  wire [15:0] _GEN_70 = 3'h0 == dstReg ? si : _GEN_62; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 46:19]
  wire [15:0] _GEN_71 = 3'h0 == dstReg ? di : _GEN_63; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 47:19]
  wire  flags_zf = result[15:0] == 16'h0; // @[src/main/scala/cpu8086/CPU8086.scala 76:21]
  wire  flags_sf = result[15]; // @[src/main/scala/cpu8086/CPU8086.scala 77:20]
  wire [1:0] _flags_pf_T_9 = result[0] + result[1]; // @[src/main/scala/cpu8086/CPU8086.scala 78:22]
  wire [1:0] _flags_pf_T_11 = result[2] + result[3]; // @[src/main/scala/cpu8086/CPU8086.scala 78:22]
  wire [2:0] _flags_pf_T_13 = _flags_pf_T_9 + _flags_pf_T_11; // @[src/main/scala/cpu8086/CPU8086.scala 78:22]
  wire [1:0] _flags_pf_T_15 = result[4] + result[5]; // @[src/main/scala/cpu8086/CPU8086.scala 78:22]
  wire [1:0] _flags_pf_T_17 = result[6] + result[7]; // @[src/main/scala/cpu8086/CPU8086.scala 78:22]
  wire [2:0] _flags_pf_T_19 = _flags_pf_T_15 + _flags_pf_T_17; // @[src/main/scala/cpu8086/CPU8086.scala 78:22]
  wire [3:0] _flags_pf_T_21 = _flags_pf_T_13 + _flags_pf_T_19; // @[src/main/scala/cpu8086/CPU8086.scala 78:22]
  wire [3:0] _GEN_261 = _flags_pf_T_21 % 4'h2; // @[src/main/scala/cpu8086/CPU8086.scala 78:37]
  wire  flags_pf = _GEN_261[1:0] == 2'h0; // @[src/main/scala/cpu8086/CPU8086.scala 78:43]
  wire [16:0] _flags_T_1 = {4'h0,overflow,4'h0,flags_sf,flags_zf,1'h0,2'h0,flags_pf,1'h0,carryOut}; // @[src/main/scala/cpu8086/CPU8086.scala 80:8]
  wire [16:0] result_1 = dst - srcVal; // @[src/main/scala/cpu8086/CPU8086.scala 220:28]
  wire  carryOut_1 = dst < srcVal; // @[src/main/scala/cpu8086/CPU8086.scala 221:30]
  wire  overflow_1 = dst[15] != srcVal[15] & dst[15] != result_1[15]; // @[src/main/scala/cpu8086/CPU8086.scala 222:48]
  wire [15:0] _GEN_72 = 3'h7 == dstReg ? result_1[15:0] : di; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 118:20 47:19]
  wire [15:0] _GEN_73 = 3'h6 == dstReg ? result_1[15:0] : si; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 117:20 46:19]
  wire [15:0] _GEN_74 = 3'h6 == dstReg ? di : _GEN_72; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 47:19]
  wire [15:0] _GEN_75 = 3'h5 == dstReg ? result_1[15:0] : bp; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 116:20 45:19]
  wire [15:0] _GEN_76 = 3'h5 == dstReg ? si : _GEN_73; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 46:19]
  wire [15:0] _GEN_77 = 3'h5 == dstReg ? di : _GEN_74; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 47:19]
  wire [15:0] _GEN_78 = 3'h4 == dstReg ? result_1[15:0] : sp; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 115:20 44:19]
  wire [15:0] _GEN_79 = 3'h4 == dstReg ? bp : _GEN_75; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 45:19]
  wire [15:0] _GEN_80 = 3'h4 == dstReg ? si : _GEN_76; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 46:19]
  wire [15:0] _GEN_81 = 3'h4 == dstReg ? di : _GEN_77; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 47:19]
  wire [15:0] _GEN_82 = 3'h3 == dstReg ? result_1[15:0] : bx; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 114:20 41:19]
  wire [15:0] _GEN_83 = 3'h3 == dstReg ? sp : _GEN_78; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 44:19]
  wire [15:0] _GEN_84 = 3'h3 == dstReg ? bp : _GEN_79; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 45:19]
  wire [15:0] _GEN_85 = 3'h3 == dstReg ? si : _GEN_80; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 46:19]
  wire [15:0] _GEN_86 = 3'h3 == dstReg ? di : _GEN_81; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 47:19]
  wire [15:0] _GEN_87 = 3'h2 == dstReg ? result_1[15:0] : dx; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 113:20 43:19]
  wire [15:0] _GEN_88 = 3'h2 == dstReg ? bx : _GEN_82; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 41:19]
  wire [15:0] _GEN_89 = 3'h2 == dstReg ? sp : _GEN_83; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 44:19]
  wire [15:0] _GEN_90 = 3'h2 == dstReg ? bp : _GEN_84; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 45:19]
  wire [15:0] _GEN_91 = 3'h2 == dstReg ? si : _GEN_85; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 46:19]
  wire [15:0] _GEN_92 = 3'h2 == dstReg ? di : _GEN_86; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 47:19]
  wire [15:0] _GEN_93 = 3'h1 == dstReg ? result_1[15:0] : cx; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 112:20 42:19]
  wire [15:0] _GEN_94 = 3'h1 == dstReg ? dx : _GEN_87; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 43:19]
  wire [15:0] _GEN_95 = 3'h1 == dstReg ? bx : _GEN_88; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 41:19]
  wire [15:0] _GEN_96 = 3'h1 == dstReg ? sp : _GEN_89; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 44:19]
  wire [15:0] _GEN_97 = 3'h1 == dstReg ? bp : _GEN_90; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 45:19]
  wire [15:0] _GEN_98 = 3'h1 == dstReg ? si : _GEN_91; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 46:19]
  wire [15:0] _GEN_99 = 3'h1 == dstReg ? di : _GEN_92; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 47:19]
  wire [15:0] _GEN_100 = 3'h0 == dstReg ? result_1[15:0] : ax; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 111:20 40:19]
  wire [15:0] _GEN_101 = 3'h0 == dstReg ? cx : _GEN_93; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 42:19]
  wire [15:0] _GEN_102 = 3'h0 == dstReg ? dx : _GEN_94; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 43:19]
  wire [15:0] _GEN_103 = 3'h0 == dstReg ? bx : _GEN_95; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 41:19]
  wire [15:0] _GEN_104 = 3'h0 == dstReg ? sp : _GEN_96; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 44:19]
  wire [15:0] _GEN_105 = 3'h0 == dstReg ? bp : _GEN_97; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 45:19]
  wire [15:0] _GEN_106 = 3'h0 == dstReg ? si : _GEN_98; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 46:19]
  wire [15:0] _GEN_107 = 3'h0 == dstReg ? di : _GEN_99; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 47:19]
  wire  flags_zf_1 = result_1[15:0] == 16'h0; // @[src/main/scala/cpu8086/CPU8086.scala 76:21]
  wire  flags_sf_1 = result_1[15]; // @[src/main/scala/cpu8086/CPU8086.scala 77:20]
  wire [1:0] _flags_pf_T_33 = result_1[0] + result_1[1]; // @[src/main/scala/cpu8086/CPU8086.scala 78:22]
  wire [1:0] _flags_pf_T_35 = result_1[2] + result_1[3]; // @[src/main/scala/cpu8086/CPU8086.scala 78:22]
  wire [2:0] _flags_pf_T_37 = _flags_pf_T_33 + _flags_pf_T_35; // @[src/main/scala/cpu8086/CPU8086.scala 78:22]
  wire [1:0] _flags_pf_T_39 = result_1[4] + result_1[5]; // @[src/main/scala/cpu8086/CPU8086.scala 78:22]
  wire [1:0] _flags_pf_T_41 = result_1[6] + result_1[7]; // @[src/main/scala/cpu8086/CPU8086.scala 78:22]
  wire [2:0] _flags_pf_T_43 = _flags_pf_T_39 + _flags_pf_T_41; // @[src/main/scala/cpu8086/CPU8086.scala 78:22]
  wire [3:0] _flags_pf_T_45 = _flags_pf_T_37 + _flags_pf_T_43; // @[src/main/scala/cpu8086/CPU8086.scala 78:22]
  wire [3:0] _GEN_268 = _flags_pf_T_45 % 4'h2; // @[src/main/scala/cpu8086/CPU8086.scala 78:37]
  wire  flags_pf_1 = _GEN_268[1:0] == 2'h0; // @[src/main/scala/cpu8086/CPU8086.scala 78:43]
  wire [16:0] _flags_T_3 = {4'h0,overflow_1,4'h0,flags_sf_1,flags_zf_1,1'h0,2'h0,flags_pf_1,1'h0,carryOut_1}; // @[src/main/scala/cpu8086/CPU8086.scala 80:8]
  wire [15:0] _ax_T_2 = ax + 16'h1; // @[src/main/scala/cpu8086/CPU8086.scala 230:31]
  wire  flags_zf_2 = _ax_T_2 == 16'h0; // @[src/main/scala/cpu8086/CPU8086.scala 76:21]
  wire  flags_sf_2 = _ax_T_2[15]; // @[src/main/scala/cpu8086/CPU8086.scala 77:20]
  wire [1:0] _flags_pf_T_57 = _ax_T_2[0] + _ax_T_2[1]; // @[src/main/scala/cpu8086/CPU8086.scala 78:22]
  wire [1:0] _flags_pf_T_59 = _ax_T_2[2] + _ax_T_2[3]; // @[src/main/scala/cpu8086/CPU8086.scala 78:22]
  wire [2:0] _flags_pf_T_61 = _flags_pf_T_57 + _flags_pf_T_59; // @[src/main/scala/cpu8086/CPU8086.scala 78:22]
  wire [1:0] _flags_pf_T_63 = _ax_T_2[4] + _ax_T_2[5]; // @[src/main/scala/cpu8086/CPU8086.scala 78:22]
  wire [1:0] _flags_pf_T_65 = _ax_T_2[6] + _ax_T_2[7]; // @[src/main/scala/cpu8086/CPU8086.scala 78:22]
  wire [2:0] _flags_pf_T_67 = _flags_pf_T_63 + _flags_pf_T_65; // @[src/main/scala/cpu8086/CPU8086.scala 78:22]
  wire [3:0] _flags_pf_T_69 = _flags_pf_T_61 + _flags_pf_T_67; // @[src/main/scala/cpu8086/CPU8086.scala 78:22]
  wire [3:0] _GEN_273 = _flags_pf_T_69 % 4'h2; // @[src/main/scala/cpu8086/CPU8086.scala 78:37]
  wire  flags_pf_2 = _GEN_273[1:0] == 2'h0; // @[src/main/scala/cpu8086/CPU8086.scala 78:43]
  wire [16:0] _flags_T_7 = {9'h0,flags_sf_2,flags_zf_2,1'h0,2'h0,flags_pf_2,1'h0,flags[0]}; // @[src/main/scala/cpu8086/CPU8086.scala 80:8]
  wire [15:0] _cx_T_2 = cx + 16'h1; // @[src/main/scala/cpu8086/CPU8086.scala 231:31]
  wire  flags_zf_3 = _cx_T_2 == 16'h0; // @[src/main/scala/cpu8086/CPU8086.scala 76:21]
  wire  flags_sf_3 = _cx_T_2[15]; // @[src/main/scala/cpu8086/CPU8086.scala 77:20]
  wire [1:0] _flags_pf_T_81 = _cx_T_2[0] + _cx_T_2[1]; // @[src/main/scala/cpu8086/CPU8086.scala 78:22]
  wire [1:0] _flags_pf_T_83 = _cx_T_2[2] + _cx_T_2[3]; // @[src/main/scala/cpu8086/CPU8086.scala 78:22]
  wire [2:0] _flags_pf_T_85 = _flags_pf_T_81 + _flags_pf_T_83; // @[src/main/scala/cpu8086/CPU8086.scala 78:22]
  wire [1:0] _flags_pf_T_87 = _cx_T_2[4] + _cx_T_2[5]; // @[src/main/scala/cpu8086/CPU8086.scala 78:22]
  wire [1:0] _flags_pf_T_89 = _cx_T_2[6] + _cx_T_2[7]; // @[src/main/scala/cpu8086/CPU8086.scala 78:22]
  wire [2:0] _flags_pf_T_91 = _flags_pf_T_87 + _flags_pf_T_89; // @[src/main/scala/cpu8086/CPU8086.scala 78:22]
  wire [3:0] _flags_pf_T_93 = _flags_pf_T_85 + _flags_pf_T_91; // @[src/main/scala/cpu8086/CPU8086.scala 78:22]
  wire [3:0] _GEN_278 = _flags_pf_T_93 % 4'h2; // @[src/main/scala/cpu8086/CPU8086.scala 78:37]
  wire  flags_pf_3 = _GEN_278[1:0] == 2'h0; // @[src/main/scala/cpu8086/CPU8086.scala 78:43]
  wire [16:0] _flags_T_11 = {9'h0,flags_sf_3,flags_zf_3,1'h0,2'h0,flags_pf_3,1'h0,flags[0]}; // @[src/main/scala/cpu8086/CPU8086.scala 80:8]
  wire [15:0] _dx_T_2 = dx + 16'h1; // @[src/main/scala/cpu8086/CPU8086.scala 232:31]
  wire  flags_zf_4 = _dx_T_2 == 16'h0; // @[src/main/scala/cpu8086/CPU8086.scala 76:21]
  wire  flags_sf_4 = _dx_T_2[15]; // @[src/main/scala/cpu8086/CPU8086.scala 77:20]
  wire [1:0] _flags_pf_T_105 = _dx_T_2[0] + _dx_T_2[1]; // @[src/main/scala/cpu8086/CPU8086.scala 78:22]
  wire [1:0] _flags_pf_T_107 = _dx_T_2[2] + _dx_T_2[3]; // @[src/main/scala/cpu8086/CPU8086.scala 78:22]
  wire [2:0] _flags_pf_T_109 = _flags_pf_T_105 + _flags_pf_T_107; // @[src/main/scala/cpu8086/CPU8086.scala 78:22]
  wire [1:0] _flags_pf_T_111 = _dx_T_2[4] + _dx_T_2[5]; // @[src/main/scala/cpu8086/CPU8086.scala 78:22]
  wire [1:0] _flags_pf_T_113 = _dx_T_2[6] + _dx_T_2[7]; // @[src/main/scala/cpu8086/CPU8086.scala 78:22]
  wire [2:0] _flags_pf_T_115 = _flags_pf_T_111 + _flags_pf_T_113; // @[src/main/scala/cpu8086/CPU8086.scala 78:22]
  wire [3:0] _flags_pf_T_117 = _flags_pf_T_109 + _flags_pf_T_115; // @[src/main/scala/cpu8086/CPU8086.scala 78:22]
  wire [3:0] _GEN_283 = _flags_pf_T_117 % 4'h2; // @[src/main/scala/cpu8086/CPU8086.scala 78:37]
  wire  flags_pf_4 = _GEN_283[1:0] == 2'h0; // @[src/main/scala/cpu8086/CPU8086.scala 78:43]
  wire [16:0] _flags_T_15 = {9'h0,flags_sf_4,flags_zf_4,1'h0,2'h0,flags_pf_4,1'h0,flags[0]}; // @[src/main/scala/cpu8086/CPU8086.scala 80:8]
  wire [15:0] _bx_T_2 = bx + 16'h1; // @[src/main/scala/cpu8086/CPU8086.scala 233:31]
  wire  flags_zf_5 = _bx_T_2 == 16'h0; // @[src/main/scala/cpu8086/CPU8086.scala 76:21]
  wire  flags_sf_5 = _bx_T_2[15]; // @[src/main/scala/cpu8086/CPU8086.scala 77:20]
  wire [1:0] _flags_pf_T_129 = _bx_T_2[0] + _bx_T_2[1]; // @[src/main/scala/cpu8086/CPU8086.scala 78:22]
  wire [1:0] _flags_pf_T_131 = _bx_T_2[2] + _bx_T_2[3]; // @[src/main/scala/cpu8086/CPU8086.scala 78:22]
  wire [2:0] _flags_pf_T_133 = _flags_pf_T_129 + _flags_pf_T_131; // @[src/main/scala/cpu8086/CPU8086.scala 78:22]
  wire [1:0] _flags_pf_T_135 = _bx_T_2[4] + _bx_T_2[5]; // @[src/main/scala/cpu8086/CPU8086.scala 78:22]
  wire [1:0] _flags_pf_T_137 = _bx_T_2[6] + _bx_T_2[7]; // @[src/main/scala/cpu8086/CPU8086.scala 78:22]
  wire [2:0] _flags_pf_T_139 = _flags_pf_T_135 + _flags_pf_T_137; // @[src/main/scala/cpu8086/CPU8086.scala 78:22]
  wire [3:0] _flags_pf_T_141 = _flags_pf_T_133 + _flags_pf_T_139; // @[src/main/scala/cpu8086/CPU8086.scala 78:22]
  wire [3:0] _GEN_288 = _flags_pf_T_141 % 4'h2; // @[src/main/scala/cpu8086/CPU8086.scala 78:37]
  wire  flags_pf_5 = _GEN_288[1:0] == 2'h0; // @[src/main/scala/cpu8086/CPU8086.scala 78:43]
  wire [16:0] _flags_T_19 = {9'h0,flags_sf_5,flags_zf_5,1'h0,2'h0,flags_pf_5,1'h0,flags[0]}; // @[src/main/scala/cpu8086/CPU8086.scala 80:8]
  wire [15:0] _sp_T_1 = sp + 16'h1; // @[src/main/scala/cpu8086/CPU8086.scala 234:31]
  wire  flags_zf_6 = _sp_T_1 == 16'h0; // @[src/main/scala/cpu8086/CPU8086.scala 76:21]
  wire  flags_sf_6 = _sp_T_1[15]; // @[src/main/scala/cpu8086/CPU8086.scala 77:20]
  wire [1:0] _flags_pf_T_153 = _sp_T_1[0] + _sp_T_1[1]; // @[src/main/scala/cpu8086/CPU8086.scala 78:22]
  wire [1:0] _flags_pf_T_155 = _sp_T_1[2] + _sp_T_1[3]; // @[src/main/scala/cpu8086/CPU8086.scala 78:22]
  wire [2:0] _flags_pf_T_157 = _flags_pf_T_153 + _flags_pf_T_155; // @[src/main/scala/cpu8086/CPU8086.scala 78:22]
  wire [1:0] _flags_pf_T_159 = _sp_T_1[4] + _sp_T_1[5]; // @[src/main/scala/cpu8086/CPU8086.scala 78:22]
  wire [1:0] _flags_pf_T_161 = _sp_T_1[6] + _sp_T_1[7]; // @[src/main/scala/cpu8086/CPU8086.scala 78:22]
  wire [2:0] _flags_pf_T_163 = _flags_pf_T_159 + _flags_pf_T_161; // @[src/main/scala/cpu8086/CPU8086.scala 78:22]
  wire [3:0] _flags_pf_T_165 = _flags_pf_T_157 + _flags_pf_T_163; // @[src/main/scala/cpu8086/CPU8086.scala 78:22]
  wire [3:0] _GEN_293 = _flags_pf_T_165 % 4'h2; // @[src/main/scala/cpu8086/CPU8086.scala 78:37]
  wire  flags_pf_6 = _GEN_293[1:0] == 2'h0; // @[src/main/scala/cpu8086/CPU8086.scala 78:43]
  wire [16:0] _flags_T_23 = {9'h0,flags_sf_6,flags_zf_6,1'h0,2'h0,flags_pf_6,1'h0,flags[0]}; // @[src/main/scala/cpu8086/CPU8086.scala 80:8]
  wire [15:0] _bp_T_1 = bp + 16'h1; // @[src/main/scala/cpu8086/CPU8086.scala 235:31]
  wire  flags_zf_7 = _bp_T_1 == 16'h0; // @[src/main/scala/cpu8086/CPU8086.scala 76:21]
  wire  flags_sf_7 = _bp_T_1[15]; // @[src/main/scala/cpu8086/CPU8086.scala 77:20]
  wire [1:0] _flags_pf_T_177 = _bp_T_1[0] + _bp_T_1[1]; // @[src/main/scala/cpu8086/CPU8086.scala 78:22]
  wire [1:0] _flags_pf_T_179 = _bp_T_1[2] + _bp_T_1[3]; // @[src/main/scala/cpu8086/CPU8086.scala 78:22]
  wire [2:0] _flags_pf_T_181 = _flags_pf_T_177 + _flags_pf_T_179; // @[src/main/scala/cpu8086/CPU8086.scala 78:22]
  wire [1:0] _flags_pf_T_183 = _bp_T_1[4] + _bp_T_1[5]; // @[src/main/scala/cpu8086/CPU8086.scala 78:22]
  wire [1:0] _flags_pf_T_185 = _bp_T_1[6] + _bp_T_1[7]; // @[src/main/scala/cpu8086/CPU8086.scala 78:22]
  wire [2:0] _flags_pf_T_187 = _flags_pf_T_183 + _flags_pf_T_185; // @[src/main/scala/cpu8086/CPU8086.scala 78:22]
  wire [3:0] _flags_pf_T_189 = _flags_pf_T_181 + _flags_pf_T_187; // @[src/main/scala/cpu8086/CPU8086.scala 78:22]
  wire [3:0] _GEN_298 = _flags_pf_T_189 % 4'h2; // @[src/main/scala/cpu8086/CPU8086.scala 78:37]
  wire  flags_pf_7 = _GEN_298[1:0] == 2'h0; // @[src/main/scala/cpu8086/CPU8086.scala 78:43]
  wire [16:0] _flags_T_27 = {9'h0,flags_sf_7,flags_zf_7,1'h0,2'h0,flags_pf_7,1'h0,flags[0]}; // @[src/main/scala/cpu8086/CPU8086.scala 80:8]
  wire [15:0] _si_T_1 = si + 16'h1; // @[src/main/scala/cpu8086/CPU8086.scala 236:31]
  wire  flags_zf_8 = _si_T_1 == 16'h0; // @[src/main/scala/cpu8086/CPU8086.scala 76:21]
  wire  flags_sf_8 = _si_T_1[15]; // @[src/main/scala/cpu8086/CPU8086.scala 77:20]
  wire [1:0] _flags_pf_T_201 = _si_T_1[0] + _si_T_1[1]; // @[src/main/scala/cpu8086/CPU8086.scala 78:22]
  wire [1:0] _flags_pf_T_203 = _si_T_1[2] + _si_T_1[3]; // @[src/main/scala/cpu8086/CPU8086.scala 78:22]
  wire [2:0] _flags_pf_T_205 = _flags_pf_T_201 + _flags_pf_T_203; // @[src/main/scala/cpu8086/CPU8086.scala 78:22]
  wire [1:0] _flags_pf_T_207 = _si_T_1[4] + _si_T_1[5]; // @[src/main/scala/cpu8086/CPU8086.scala 78:22]
  wire [1:0] _flags_pf_T_209 = _si_T_1[6] + _si_T_1[7]; // @[src/main/scala/cpu8086/CPU8086.scala 78:22]
  wire [2:0] _flags_pf_T_211 = _flags_pf_T_207 + _flags_pf_T_209; // @[src/main/scala/cpu8086/CPU8086.scala 78:22]
  wire [3:0] _flags_pf_T_213 = _flags_pf_T_205 + _flags_pf_T_211; // @[src/main/scala/cpu8086/CPU8086.scala 78:22]
  wire [3:0] _GEN_303 = _flags_pf_T_213 % 4'h2; // @[src/main/scala/cpu8086/CPU8086.scala 78:37]
  wire  flags_pf_8 = _GEN_303[1:0] == 2'h0; // @[src/main/scala/cpu8086/CPU8086.scala 78:43]
  wire [16:0] _flags_T_31 = {9'h0,flags_sf_8,flags_zf_8,1'h0,2'h0,flags_pf_8,1'h0,flags[0]}; // @[src/main/scala/cpu8086/CPU8086.scala 80:8]
  wire [15:0] _di_T_1 = di + 16'h1; // @[src/main/scala/cpu8086/CPU8086.scala 237:31]
  wire  flags_zf_9 = _di_T_1 == 16'h0; // @[src/main/scala/cpu8086/CPU8086.scala 76:21]
  wire  flags_sf_9 = _di_T_1[15]; // @[src/main/scala/cpu8086/CPU8086.scala 77:20]
  wire [1:0] _flags_pf_T_225 = _di_T_1[0] + _di_T_1[1]; // @[src/main/scala/cpu8086/CPU8086.scala 78:22]
  wire [1:0] _flags_pf_T_227 = _di_T_1[2] + _di_T_1[3]; // @[src/main/scala/cpu8086/CPU8086.scala 78:22]
  wire [2:0] _flags_pf_T_229 = _flags_pf_T_225 + _flags_pf_T_227; // @[src/main/scala/cpu8086/CPU8086.scala 78:22]
  wire [1:0] _flags_pf_T_231 = _di_T_1[4] + _di_T_1[5]; // @[src/main/scala/cpu8086/CPU8086.scala 78:22]
  wire [1:0] _flags_pf_T_233 = _di_T_1[6] + _di_T_1[7]; // @[src/main/scala/cpu8086/CPU8086.scala 78:22]
  wire [2:0] _flags_pf_T_235 = _flags_pf_T_231 + _flags_pf_T_233; // @[src/main/scala/cpu8086/CPU8086.scala 78:22]
  wire [3:0] _flags_pf_T_237 = _flags_pf_T_229 + _flags_pf_T_235; // @[src/main/scala/cpu8086/CPU8086.scala 78:22]
  wire [3:0] _GEN_308 = _flags_pf_T_237 % 4'h2; // @[src/main/scala/cpu8086/CPU8086.scala 78:37]
  wire  flags_pf_9 = _GEN_308[1:0] == 2'h0; // @[src/main/scala/cpu8086/CPU8086.scala 78:43]
  wire [16:0] _flags_T_35 = {9'h0,flags_sf_9,flags_zf_9,1'h0,2'h0,flags_pf_9,1'h0,flags[0]}; // @[src/main/scala/cpu8086/CPU8086.scala 80:8]
  wire [15:0] _ax_T_4 = ax - 16'h1; // @[src/main/scala/cpu8086/CPU8086.scala 240:31]
  wire  flags_zf_10 = _ax_T_4 == 16'h0; // @[src/main/scala/cpu8086/CPU8086.scala 76:21]
  wire  flags_sf_10 = _ax_T_4[15]; // @[src/main/scala/cpu8086/CPU8086.scala 77:20]
  wire [1:0] _flags_pf_T_249 = _ax_T_4[0] + _ax_T_4[1]; // @[src/main/scala/cpu8086/CPU8086.scala 78:22]
  wire [1:0] _flags_pf_T_251 = _ax_T_4[2] + _ax_T_4[3]; // @[src/main/scala/cpu8086/CPU8086.scala 78:22]
  wire [2:0] _flags_pf_T_253 = _flags_pf_T_249 + _flags_pf_T_251; // @[src/main/scala/cpu8086/CPU8086.scala 78:22]
  wire [1:0] _flags_pf_T_255 = _ax_T_4[4] + _ax_T_4[5]; // @[src/main/scala/cpu8086/CPU8086.scala 78:22]
  wire [1:0] _flags_pf_T_257 = _ax_T_4[6] + _ax_T_4[7]; // @[src/main/scala/cpu8086/CPU8086.scala 78:22]
  wire [2:0] _flags_pf_T_259 = _flags_pf_T_255 + _flags_pf_T_257; // @[src/main/scala/cpu8086/CPU8086.scala 78:22]
  wire [3:0] _flags_pf_T_261 = _flags_pf_T_253 + _flags_pf_T_259; // @[src/main/scala/cpu8086/CPU8086.scala 78:22]
  wire [3:0] _GEN_313 = _flags_pf_T_261 % 4'h2; // @[src/main/scala/cpu8086/CPU8086.scala 78:37]
  wire  flags_pf_10 = _GEN_313[1:0] == 2'h0; // @[src/main/scala/cpu8086/CPU8086.scala 78:43]
  wire [16:0] _flags_T_39 = {9'h0,flags_sf_10,flags_zf_10,1'h0,2'h0,flags_pf_10,1'h0,flags[0]}; // @[src/main/scala/cpu8086/CPU8086.scala 80:8]
  wire [15:0] _cx_T_4 = cx - 16'h1; // @[src/main/scala/cpu8086/CPU8086.scala 241:31]
  wire  flags_zf_11 = _cx_T_4 == 16'h0; // @[src/main/scala/cpu8086/CPU8086.scala 76:21]
  wire  flags_sf_11 = _cx_T_4[15]; // @[src/main/scala/cpu8086/CPU8086.scala 77:20]
  wire [1:0] _flags_pf_T_273 = _cx_T_4[0] + _cx_T_4[1]; // @[src/main/scala/cpu8086/CPU8086.scala 78:22]
  wire [1:0] _flags_pf_T_275 = _cx_T_4[2] + _cx_T_4[3]; // @[src/main/scala/cpu8086/CPU8086.scala 78:22]
  wire [2:0] _flags_pf_T_277 = _flags_pf_T_273 + _flags_pf_T_275; // @[src/main/scala/cpu8086/CPU8086.scala 78:22]
  wire [1:0] _flags_pf_T_279 = _cx_T_4[4] + _cx_T_4[5]; // @[src/main/scala/cpu8086/CPU8086.scala 78:22]
  wire [1:0] _flags_pf_T_281 = _cx_T_4[6] + _cx_T_4[7]; // @[src/main/scala/cpu8086/CPU8086.scala 78:22]
  wire [2:0] _flags_pf_T_283 = _flags_pf_T_279 + _flags_pf_T_281; // @[src/main/scala/cpu8086/CPU8086.scala 78:22]
  wire [3:0] _flags_pf_T_285 = _flags_pf_T_277 + _flags_pf_T_283; // @[src/main/scala/cpu8086/CPU8086.scala 78:22]
  wire [3:0] _GEN_318 = _flags_pf_T_285 % 4'h2; // @[src/main/scala/cpu8086/CPU8086.scala 78:37]
  wire  flags_pf_11 = _GEN_318[1:0] == 2'h0; // @[src/main/scala/cpu8086/CPU8086.scala 78:43]
  wire [16:0] _flags_T_43 = {9'h0,flags_sf_11,flags_zf_11,1'h0,2'h0,flags_pf_11,1'h0,flags[0]}; // @[src/main/scala/cpu8086/CPU8086.scala 80:8]
  wire [15:0] _dx_T_4 = dx - 16'h1; // @[src/main/scala/cpu8086/CPU8086.scala 242:31]
  wire  flags_zf_12 = _dx_T_4 == 16'h0; // @[src/main/scala/cpu8086/CPU8086.scala 76:21]
  wire  flags_sf_12 = _dx_T_4[15]; // @[src/main/scala/cpu8086/CPU8086.scala 77:20]
  wire [1:0] _flags_pf_T_297 = _dx_T_4[0] + _dx_T_4[1]; // @[src/main/scala/cpu8086/CPU8086.scala 78:22]
  wire [1:0] _flags_pf_T_299 = _dx_T_4[2] + _dx_T_4[3]; // @[src/main/scala/cpu8086/CPU8086.scala 78:22]
  wire [2:0] _flags_pf_T_301 = _flags_pf_T_297 + _flags_pf_T_299; // @[src/main/scala/cpu8086/CPU8086.scala 78:22]
  wire [1:0] _flags_pf_T_303 = _dx_T_4[4] + _dx_T_4[5]; // @[src/main/scala/cpu8086/CPU8086.scala 78:22]
  wire [1:0] _flags_pf_T_305 = _dx_T_4[6] + _dx_T_4[7]; // @[src/main/scala/cpu8086/CPU8086.scala 78:22]
  wire [2:0] _flags_pf_T_307 = _flags_pf_T_303 + _flags_pf_T_305; // @[src/main/scala/cpu8086/CPU8086.scala 78:22]
  wire [3:0] _flags_pf_T_309 = _flags_pf_T_301 + _flags_pf_T_307; // @[src/main/scala/cpu8086/CPU8086.scala 78:22]
  wire [3:0] _GEN_325 = _flags_pf_T_309 % 4'h2; // @[src/main/scala/cpu8086/CPU8086.scala 78:37]
  wire  flags_pf_12 = _GEN_325[1:0] == 2'h0; // @[src/main/scala/cpu8086/CPU8086.scala 78:43]
  wire [16:0] _flags_T_47 = {9'h0,flags_sf_12,flags_zf_12,1'h0,2'h0,flags_pf_12,1'h0,flags[0]}; // @[src/main/scala/cpu8086/CPU8086.scala 80:8]
  wire [15:0] _bx_T_4 = bx - 16'h1; // @[src/main/scala/cpu8086/CPU8086.scala 243:31]
  wire  flags_zf_13 = _bx_T_4 == 16'h0; // @[src/main/scala/cpu8086/CPU8086.scala 76:21]
  wire  flags_sf_13 = _bx_T_4[15]; // @[src/main/scala/cpu8086/CPU8086.scala 77:20]
  wire [1:0] _flags_pf_T_321 = _bx_T_4[0] + _bx_T_4[1]; // @[src/main/scala/cpu8086/CPU8086.scala 78:22]
  wire [1:0] _flags_pf_T_323 = _bx_T_4[2] + _bx_T_4[3]; // @[src/main/scala/cpu8086/CPU8086.scala 78:22]
  wire [2:0] _flags_pf_T_325 = _flags_pf_T_321 + _flags_pf_T_323; // @[src/main/scala/cpu8086/CPU8086.scala 78:22]
  wire [1:0] _flags_pf_T_327 = _bx_T_4[4] + _bx_T_4[5]; // @[src/main/scala/cpu8086/CPU8086.scala 78:22]
  wire [1:0] _flags_pf_T_329 = _bx_T_4[6] + _bx_T_4[7]; // @[src/main/scala/cpu8086/CPU8086.scala 78:22]
  wire [2:0] _flags_pf_T_331 = _flags_pf_T_327 + _flags_pf_T_329; // @[src/main/scala/cpu8086/CPU8086.scala 78:22]
  wire [3:0] _flags_pf_T_333 = _flags_pf_T_325 + _flags_pf_T_331; // @[src/main/scala/cpu8086/CPU8086.scala 78:22]
  wire [3:0] _GEN_330 = _flags_pf_T_333 % 4'h2; // @[src/main/scala/cpu8086/CPU8086.scala 78:37]
  wire  flags_pf_13 = _GEN_330[1:0] == 2'h0; // @[src/main/scala/cpu8086/CPU8086.scala 78:43]
  wire [16:0] _flags_T_51 = {9'h0,flags_sf_13,flags_zf_13,1'h0,2'h0,flags_pf_13,1'h0,flags[0]}; // @[src/main/scala/cpu8086/CPU8086.scala 80:8]
  wire [15:0] _sp_T_3 = sp - 16'h1; // @[src/main/scala/cpu8086/CPU8086.scala 244:31]
  wire  flags_zf_14 = _sp_T_3 == 16'h0; // @[src/main/scala/cpu8086/CPU8086.scala 76:21]
  wire  flags_sf_14 = _sp_T_3[15]; // @[src/main/scala/cpu8086/CPU8086.scala 77:20]
  wire [1:0] _flags_pf_T_345 = _sp_T_3[0] + _sp_T_3[1]; // @[src/main/scala/cpu8086/CPU8086.scala 78:22]
  wire [1:0] _flags_pf_T_347 = _sp_T_3[2] + _sp_T_3[3]; // @[src/main/scala/cpu8086/CPU8086.scala 78:22]
  wire [2:0] _flags_pf_T_349 = _flags_pf_T_345 + _flags_pf_T_347; // @[src/main/scala/cpu8086/CPU8086.scala 78:22]
  wire [1:0] _flags_pf_T_351 = _sp_T_3[4] + _sp_T_3[5]; // @[src/main/scala/cpu8086/CPU8086.scala 78:22]
  wire [1:0] _flags_pf_T_353 = _sp_T_3[6] + _sp_T_3[7]; // @[src/main/scala/cpu8086/CPU8086.scala 78:22]
  wire [2:0] _flags_pf_T_355 = _flags_pf_T_351 + _flags_pf_T_353; // @[src/main/scala/cpu8086/CPU8086.scala 78:22]
  wire [3:0] _flags_pf_T_357 = _flags_pf_T_349 + _flags_pf_T_355; // @[src/main/scala/cpu8086/CPU8086.scala 78:22]
  wire [3:0] _GEN_335 = _flags_pf_T_357 % 4'h2; // @[src/main/scala/cpu8086/CPU8086.scala 78:37]
  wire  flags_pf_14 = _GEN_335[1:0] == 2'h0; // @[src/main/scala/cpu8086/CPU8086.scala 78:43]
  wire [16:0] _flags_T_55 = {9'h0,flags_sf_14,flags_zf_14,1'h0,2'h0,flags_pf_14,1'h0,flags[0]}; // @[src/main/scala/cpu8086/CPU8086.scala 80:8]
  wire [15:0] _bp_T_3 = bp - 16'h1; // @[src/main/scala/cpu8086/CPU8086.scala 245:31]
  wire  flags_zf_15 = _bp_T_3 == 16'h0; // @[src/main/scala/cpu8086/CPU8086.scala 76:21]
  wire  flags_sf_15 = _bp_T_3[15]; // @[src/main/scala/cpu8086/CPU8086.scala 77:20]
  wire [1:0] _flags_pf_T_369 = _bp_T_3[0] + _bp_T_3[1]; // @[src/main/scala/cpu8086/CPU8086.scala 78:22]
  wire [1:0] _flags_pf_T_371 = _bp_T_3[2] + _bp_T_3[3]; // @[src/main/scala/cpu8086/CPU8086.scala 78:22]
  wire [2:0] _flags_pf_T_373 = _flags_pf_T_369 + _flags_pf_T_371; // @[src/main/scala/cpu8086/CPU8086.scala 78:22]
  wire [1:0] _flags_pf_T_375 = _bp_T_3[4] + _bp_T_3[5]; // @[src/main/scala/cpu8086/CPU8086.scala 78:22]
  wire [1:0] _flags_pf_T_377 = _bp_T_3[6] + _bp_T_3[7]; // @[src/main/scala/cpu8086/CPU8086.scala 78:22]
  wire [2:0] _flags_pf_T_379 = _flags_pf_T_375 + _flags_pf_T_377; // @[src/main/scala/cpu8086/CPU8086.scala 78:22]
  wire [3:0] _flags_pf_T_381 = _flags_pf_T_373 + _flags_pf_T_379; // @[src/main/scala/cpu8086/CPU8086.scala 78:22]
  wire [3:0] _GEN_340 = _flags_pf_T_381 % 4'h2; // @[src/main/scala/cpu8086/CPU8086.scala 78:37]
  wire  flags_pf_15 = _GEN_340[1:0] == 2'h0; // @[src/main/scala/cpu8086/CPU8086.scala 78:43]
  wire [16:0] _flags_T_59 = {9'h0,flags_sf_15,flags_zf_15,1'h0,2'h0,flags_pf_15,1'h0,flags[0]}; // @[src/main/scala/cpu8086/CPU8086.scala 80:8]
  wire [15:0] _si_T_3 = si - 16'h1; // @[src/main/scala/cpu8086/CPU8086.scala 246:31]
  wire  flags_zf_16 = _si_T_3 == 16'h0; // @[src/main/scala/cpu8086/CPU8086.scala 76:21]
  wire  flags_sf_16 = _si_T_3[15]; // @[src/main/scala/cpu8086/CPU8086.scala 77:20]
  wire [1:0] _flags_pf_T_393 = _si_T_3[0] + _si_T_3[1]; // @[src/main/scala/cpu8086/CPU8086.scala 78:22]
  wire [1:0] _flags_pf_T_395 = _si_T_3[2] + _si_T_3[3]; // @[src/main/scala/cpu8086/CPU8086.scala 78:22]
  wire [2:0] _flags_pf_T_397 = _flags_pf_T_393 + _flags_pf_T_395; // @[src/main/scala/cpu8086/CPU8086.scala 78:22]
  wire [1:0] _flags_pf_T_399 = _si_T_3[4] + _si_T_3[5]; // @[src/main/scala/cpu8086/CPU8086.scala 78:22]
  wire [1:0] _flags_pf_T_401 = _si_T_3[6] + _si_T_3[7]; // @[src/main/scala/cpu8086/CPU8086.scala 78:22]
  wire [2:0] _flags_pf_T_403 = _flags_pf_T_399 + _flags_pf_T_401; // @[src/main/scala/cpu8086/CPU8086.scala 78:22]
  wire [3:0] _flags_pf_T_405 = _flags_pf_T_397 + _flags_pf_T_403; // @[src/main/scala/cpu8086/CPU8086.scala 78:22]
  wire [3:0] _GEN_346 = _flags_pf_T_405 % 4'h2; // @[src/main/scala/cpu8086/CPU8086.scala 78:37]
  wire  flags_pf_16 = _GEN_346[1:0] == 2'h0; // @[src/main/scala/cpu8086/CPU8086.scala 78:43]
  wire [16:0] _flags_T_63 = {9'h0,flags_sf_16,flags_zf_16,1'h0,2'h0,flags_pf_16,1'h0,flags[0]}; // @[src/main/scala/cpu8086/CPU8086.scala 80:8]
  wire [15:0] _di_T_3 = di - 16'h1; // @[src/main/scala/cpu8086/CPU8086.scala 247:31]
  wire  flags_zf_17 = _di_T_3 == 16'h0; // @[src/main/scala/cpu8086/CPU8086.scala 76:21]
  wire  flags_sf_17 = _di_T_3[15]; // @[src/main/scala/cpu8086/CPU8086.scala 77:20]
  wire [1:0] _flags_pf_T_417 = _di_T_3[0] + _di_T_3[1]; // @[src/main/scala/cpu8086/CPU8086.scala 78:22]
  wire [1:0] _flags_pf_T_419 = _di_T_3[2] + _di_T_3[3]; // @[src/main/scala/cpu8086/CPU8086.scala 78:22]
  wire [2:0] _flags_pf_T_421 = _flags_pf_T_417 + _flags_pf_T_419; // @[src/main/scala/cpu8086/CPU8086.scala 78:22]
  wire [1:0] _flags_pf_T_423 = _di_T_3[4] + _di_T_3[5]; // @[src/main/scala/cpu8086/CPU8086.scala 78:22]
  wire [1:0] _flags_pf_T_425 = _di_T_3[6] + _di_T_3[7]; // @[src/main/scala/cpu8086/CPU8086.scala 78:22]
  wire [2:0] _flags_pf_T_427 = _flags_pf_T_423 + _flags_pf_T_425; // @[src/main/scala/cpu8086/CPU8086.scala 78:22]
  wire [3:0] _flags_pf_T_429 = _flags_pf_T_421 + _flags_pf_T_427; // @[src/main/scala/cpu8086/CPU8086.scala 78:22]
  wire [3:0] _GEN_359 = _flags_pf_T_429 % 4'h2; // @[src/main/scala/cpu8086/CPU8086.scala 78:37]
  wire  flags_pf_17 = _GEN_359[1:0] == 2'h0; // @[src/main/scala/cpu8086/CPU8086.scala 78:43]
  wire [16:0] _flags_T_67 = {9'h0,flags_sf_17,flags_zf_17,1'h0,2'h0,flags_pf_17,1'h0,flags[0]}; // @[src/main/scala/cpu8086/CPU8086.scala 80:8]
  wire [15:0] result_3 = dst & srcVal; // @[src/main/scala/cpu8086/CPU8086.scala 267:28]
  wire [15:0] _GEN_108 = 3'h7 == dstReg ? result_3 : di; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 118:20 47:19]
  wire [15:0] _GEN_109 = 3'h6 == dstReg ? result_3 : si; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 117:20 46:19]
  wire [15:0] _GEN_110 = 3'h6 == dstReg ? di : _GEN_108; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 47:19]
  wire [15:0] _GEN_111 = 3'h5 == dstReg ? result_3 : bp; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 116:20 45:19]
  wire [15:0] _GEN_112 = 3'h5 == dstReg ? si : _GEN_109; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 46:19]
  wire [15:0] _GEN_113 = 3'h5 == dstReg ? di : _GEN_110; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 47:19]
  wire [15:0] _GEN_114 = 3'h4 == dstReg ? result_3 : sp; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 115:20 44:19]
  wire [15:0] _GEN_115 = 3'h4 == dstReg ? bp : _GEN_111; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 45:19]
  wire [15:0] _GEN_116 = 3'h4 == dstReg ? si : _GEN_112; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 46:19]
  wire [15:0] _GEN_117 = 3'h4 == dstReg ? di : _GEN_113; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 47:19]
  wire [15:0] _GEN_118 = 3'h3 == dstReg ? result_3 : bx; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 114:20 41:19]
  wire [15:0] _GEN_119 = 3'h3 == dstReg ? sp : _GEN_114; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 44:19]
  wire [15:0] _GEN_120 = 3'h3 == dstReg ? bp : _GEN_115; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 45:19]
  wire [15:0] _GEN_121 = 3'h3 == dstReg ? si : _GEN_116; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 46:19]
  wire [15:0] _GEN_122 = 3'h3 == dstReg ? di : _GEN_117; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 47:19]
  wire [15:0] _GEN_123 = 3'h2 == dstReg ? result_3 : dx; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 113:20 43:19]
  wire [15:0] _GEN_124 = 3'h2 == dstReg ? bx : _GEN_118; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 41:19]
  wire [15:0] _GEN_125 = 3'h2 == dstReg ? sp : _GEN_119; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 44:19]
  wire [15:0] _GEN_126 = 3'h2 == dstReg ? bp : _GEN_120; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 45:19]
  wire [15:0] _GEN_127 = 3'h2 == dstReg ? si : _GEN_121; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 46:19]
  wire [15:0] _GEN_128 = 3'h2 == dstReg ? di : _GEN_122; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 47:19]
  wire [15:0] _GEN_129 = 3'h1 == dstReg ? result_3 : cx; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 112:20 42:19]
  wire [15:0] _GEN_130 = 3'h1 == dstReg ? dx : _GEN_123; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 43:19]
  wire [15:0] _GEN_131 = 3'h1 == dstReg ? bx : _GEN_124; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 41:19]
  wire [15:0] _GEN_132 = 3'h1 == dstReg ? sp : _GEN_125; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 44:19]
  wire [15:0] _GEN_133 = 3'h1 == dstReg ? bp : _GEN_126; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 45:19]
  wire [15:0] _GEN_134 = 3'h1 == dstReg ? si : _GEN_127; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 46:19]
  wire [15:0] _GEN_135 = 3'h1 == dstReg ? di : _GEN_128; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 47:19]
  wire [15:0] _GEN_136 = 3'h0 == dstReg ? result_3 : ax; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 111:20 40:19]
  wire [15:0] _GEN_137 = 3'h0 == dstReg ? cx : _GEN_129; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 42:19]
  wire [15:0] _GEN_138 = 3'h0 == dstReg ? dx : _GEN_130; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 43:19]
  wire [15:0] _GEN_139 = 3'h0 == dstReg ? bx : _GEN_131; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 41:19]
  wire [15:0] _GEN_140 = 3'h0 == dstReg ? sp : _GEN_132; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 44:19]
  wire [15:0] _GEN_141 = 3'h0 == dstReg ? bp : _GEN_133; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 45:19]
  wire [15:0] _GEN_142 = 3'h0 == dstReg ? si : _GEN_134; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 46:19]
  wire [15:0] _GEN_143 = 3'h0 == dstReg ? di : _GEN_135; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 47:19]
  wire  flags_zf_19 = result_3 == 16'h0; // @[src/main/scala/cpu8086/CPU8086.scala 76:21]
  wire  flags_sf_19 = result_3[15]; // @[src/main/scala/cpu8086/CPU8086.scala 77:20]
  wire [1:0] _flags_pf_T_465 = result_3[0] + result_3[1]; // @[src/main/scala/cpu8086/CPU8086.scala 78:22]
  wire [1:0] _flags_pf_T_467 = result_3[2] + result_3[3]; // @[src/main/scala/cpu8086/CPU8086.scala 78:22]
  wire [2:0] _flags_pf_T_469 = _flags_pf_T_465 + _flags_pf_T_467; // @[src/main/scala/cpu8086/CPU8086.scala 78:22]
  wire [1:0] _flags_pf_T_471 = result_3[4] + result_3[5]; // @[src/main/scala/cpu8086/CPU8086.scala 78:22]
  wire [1:0] _flags_pf_T_473 = result_3[6] + result_3[7]; // @[src/main/scala/cpu8086/CPU8086.scala 78:22]
  wire [2:0] _flags_pf_T_475 = _flags_pf_T_471 + _flags_pf_T_473; // @[src/main/scala/cpu8086/CPU8086.scala 78:22]
  wire [3:0] _flags_pf_T_477 = _flags_pf_T_469 + _flags_pf_T_475; // @[src/main/scala/cpu8086/CPU8086.scala 78:22]
  wire [3:0] _GEN_372 = _flags_pf_T_477 % 4'h2; // @[src/main/scala/cpu8086/CPU8086.scala 78:37]
  wire  flags_pf_19 = _GEN_372[1:0] == 2'h0; // @[src/main/scala/cpu8086/CPU8086.scala 78:43]
  wire [16:0] _flags_T_70 = {9'h0,flags_sf_19,flags_zf_19,1'h0,2'h0,flags_pf_19,2'h0}; // @[src/main/scala/cpu8086/CPU8086.scala 80:8]
  wire [15:0] result_4 = dst | srcVal; // @[src/main/scala/cpu8086/CPU8086.scala 278:28]
  wire [15:0] _GEN_144 = 3'h7 == dstReg ? result_4 : di; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 118:20 47:19]
  wire [15:0] _GEN_145 = 3'h6 == dstReg ? result_4 : si; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 117:20 46:19]
  wire [15:0] _GEN_146 = 3'h6 == dstReg ? di : _GEN_144; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 47:19]
  wire [15:0] _GEN_147 = 3'h5 == dstReg ? result_4 : bp; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 116:20 45:19]
  wire [15:0] _GEN_148 = 3'h5 == dstReg ? si : _GEN_145; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 46:19]
  wire [15:0] _GEN_149 = 3'h5 == dstReg ? di : _GEN_146; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 47:19]
  wire [15:0] _GEN_150 = 3'h4 == dstReg ? result_4 : sp; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 115:20 44:19]
  wire [15:0] _GEN_151 = 3'h4 == dstReg ? bp : _GEN_147; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 45:19]
  wire [15:0] _GEN_152 = 3'h4 == dstReg ? si : _GEN_148; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 46:19]
  wire [15:0] _GEN_153 = 3'h4 == dstReg ? di : _GEN_149; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 47:19]
  wire [15:0] _GEN_154 = 3'h3 == dstReg ? result_4 : bx; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 114:20 41:19]
  wire [15:0] _GEN_155 = 3'h3 == dstReg ? sp : _GEN_150; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 44:19]
  wire [15:0] _GEN_156 = 3'h3 == dstReg ? bp : _GEN_151; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 45:19]
  wire [15:0] _GEN_157 = 3'h3 == dstReg ? si : _GEN_152; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 46:19]
  wire [15:0] _GEN_158 = 3'h3 == dstReg ? di : _GEN_153; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 47:19]
  wire [15:0] _GEN_159 = 3'h2 == dstReg ? result_4 : dx; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 113:20 43:19]
  wire [15:0] _GEN_160 = 3'h2 == dstReg ? bx : _GEN_154; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 41:19]
  wire [15:0] _GEN_161 = 3'h2 == dstReg ? sp : _GEN_155; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 44:19]
  wire [15:0] _GEN_162 = 3'h2 == dstReg ? bp : _GEN_156; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 45:19]
  wire [15:0] _GEN_163 = 3'h2 == dstReg ? si : _GEN_157; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 46:19]
  wire [15:0] _GEN_164 = 3'h2 == dstReg ? di : _GEN_158; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 47:19]
  wire [15:0] _GEN_165 = 3'h1 == dstReg ? result_4 : cx; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 112:20 42:19]
  wire [15:0] _GEN_166 = 3'h1 == dstReg ? dx : _GEN_159; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 43:19]
  wire [15:0] _GEN_167 = 3'h1 == dstReg ? bx : _GEN_160; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 41:19]
  wire [15:0] _GEN_168 = 3'h1 == dstReg ? sp : _GEN_161; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 44:19]
  wire [15:0] _GEN_169 = 3'h1 == dstReg ? bp : _GEN_162; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 45:19]
  wire [15:0] _GEN_170 = 3'h1 == dstReg ? si : _GEN_163; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 46:19]
  wire [15:0] _GEN_171 = 3'h1 == dstReg ? di : _GEN_164; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 47:19]
  wire [15:0] _GEN_172 = 3'h0 == dstReg ? result_4 : ax; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 111:20 40:19]
  wire [15:0] _GEN_173 = 3'h0 == dstReg ? cx : _GEN_165; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 42:19]
  wire [15:0] _GEN_174 = 3'h0 == dstReg ? dx : _GEN_166; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 43:19]
  wire [15:0] _GEN_175 = 3'h0 == dstReg ? bx : _GEN_167; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 41:19]
  wire [15:0] _GEN_176 = 3'h0 == dstReg ? sp : _GEN_168; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 44:19]
  wire [15:0] _GEN_177 = 3'h0 == dstReg ? bp : _GEN_169; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 45:19]
  wire [15:0] _GEN_178 = 3'h0 == dstReg ? si : _GEN_170; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 46:19]
  wire [15:0] _GEN_179 = 3'h0 == dstReg ? di : _GEN_171; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 47:19]
  wire  flags_zf_20 = result_4 == 16'h0; // @[src/main/scala/cpu8086/CPU8086.scala 76:21]
  wire  flags_sf_20 = result_4[15]; // @[src/main/scala/cpu8086/CPU8086.scala 77:20]
  wire [1:0] _flags_pf_T_489 = result_4[0] + result_4[1]; // @[src/main/scala/cpu8086/CPU8086.scala 78:22]
  wire [1:0] _flags_pf_T_491 = result_4[2] + result_4[3]; // @[src/main/scala/cpu8086/CPU8086.scala 78:22]
  wire [2:0] _flags_pf_T_493 = _flags_pf_T_489 + _flags_pf_T_491; // @[src/main/scala/cpu8086/CPU8086.scala 78:22]
  wire [1:0] _flags_pf_T_495 = result_4[4] + result_4[5]; // @[src/main/scala/cpu8086/CPU8086.scala 78:22]
  wire [1:0] _flags_pf_T_497 = result_4[6] + result_4[7]; // @[src/main/scala/cpu8086/CPU8086.scala 78:22]
  wire [2:0] _flags_pf_T_499 = _flags_pf_T_495 + _flags_pf_T_497; // @[src/main/scala/cpu8086/CPU8086.scala 78:22]
  wire [3:0] _flags_pf_T_501 = _flags_pf_T_493 + _flags_pf_T_499; // @[src/main/scala/cpu8086/CPU8086.scala 78:22]
  wire [3:0] _GEN_385 = _flags_pf_T_501 % 4'h2; // @[src/main/scala/cpu8086/CPU8086.scala 78:37]
  wire  flags_pf_20 = _GEN_385[1:0] == 2'h0; // @[src/main/scala/cpu8086/CPU8086.scala 78:43]
  wire [16:0] _flags_T_71 = {9'h0,flags_sf_20,flags_zf_20,1'h0,2'h0,flags_pf_20,2'h0}; // @[src/main/scala/cpu8086/CPU8086.scala 80:8]
  wire [15:0] result_5 = dst ^ srcVal; // @[src/main/scala/cpu8086/CPU8086.scala 289:28]
  wire [15:0] _GEN_180 = 3'h7 == dstReg ? result_5 : di; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 118:20 47:19]
  wire [15:0] _GEN_181 = 3'h6 == dstReg ? result_5 : si; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 117:20 46:19]
  wire [15:0] _GEN_182 = 3'h6 == dstReg ? di : _GEN_180; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 47:19]
  wire [15:0] _GEN_183 = 3'h5 == dstReg ? result_5 : bp; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 116:20 45:19]
  wire [15:0] _GEN_184 = 3'h5 == dstReg ? si : _GEN_181; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 46:19]
  wire [15:0] _GEN_185 = 3'h5 == dstReg ? di : _GEN_182; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 47:19]
  wire [15:0] _GEN_186 = 3'h4 == dstReg ? result_5 : sp; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 115:20 44:19]
  wire [15:0] _GEN_187 = 3'h4 == dstReg ? bp : _GEN_183; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 45:19]
  wire [15:0] _GEN_188 = 3'h4 == dstReg ? si : _GEN_184; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 46:19]
  wire [15:0] _GEN_189 = 3'h4 == dstReg ? di : _GEN_185; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 47:19]
  wire [15:0] _GEN_190 = 3'h3 == dstReg ? result_5 : bx; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 114:20 41:19]
  wire [15:0] _GEN_191 = 3'h3 == dstReg ? sp : _GEN_186; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 44:19]
  wire [15:0] _GEN_192 = 3'h3 == dstReg ? bp : _GEN_187; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 45:19]
  wire [15:0] _GEN_193 = 3'h3 == dstReg ? si : _GEN_188; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 46:19]
  wire [15:0] _GEN_194 = 3'h3 == dstReg ? di : _GEN_189; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 47:19]
  wire [15:0] _GEN_195 = 3'h2 == dstReg ? result_5 : dx; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 113:20 43:19]
  wire [15:0] _GEN_196 = 3'h2 == dstReg ? bx : _GEN_190; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 41:19]
  wire [15:0] _GEN_197 = 3'h2 == dstReg ? sp : _GEN_191; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 44:19]
  wire [15:0] _GEN_198 = 3'h2 == dstReg ? bp : _GEN_192; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 45:19]
  wire [15:0] _GEN_199 = 3'h2 == dstReg ? si : _GEN_193; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 46:19]
  wire [15:0] _GEN_200 = 3'h2 == dstReg ? di : _GEN_194; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 47:19]
  wire [15:0] _GEN_201 = 3'h1 == dstReg ? result_5 : cx; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 112:20 42:19]
  wire [15:0] _GEN_202 = 3'h1 == dstReg ? dx : _GEN_195; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 43:19]
  wire [15:0] _GEN_203 = 3'h1 == dstReg ? bx : _GEN_196; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 41:19]
  wire [15:0] _GEN_204 = 3'h1 == dstReg ? sp : _GEN_197; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 44:19]
  wire [15:0] _GEN_205 = 3'h1 == dstReg ? bp : _GEN_198; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 45:19]
  wire [15:0] _GEN_206 = 3'h1 == dstReg ? si : _GEN_199; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 46:19]
  wire [15:0] _GEN_207 = 3'h1 == dstReg ? di : _GEN_200; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 47:19]
  wire [15:0] _GEN_208 = 3'h0 == dstReg ? result_5 : ax; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 111:20 40:19]
  wire [15:0] _GEN_209 = 3'h0 == dstReg ? cx : _GEN_201; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 42:19]
  wire [15:0] _GEN_210 = 3'h0 == dstReg ? dx : _GEN_202; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 43:19]
  wire [15:0] _GEN_211 = 3'h0 == dstReg ? bx : _GEN_203; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 41:19]
  wire [15:0] _GEN_212 = 3'h0 == dstReg ? sp : _GEN_204; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 44:19]
  wire [15:0] _GEN_213 = 3'h0 == dstReg ? bp : _GEN_205; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 45:19]
  wire [15:0] _GEN_214 = 3'h0 == dstReg ? si : _GEN_206; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 46:19]
  wire [15:0] _GEN_215 = 3'h0 == dstReg ? di : _GEN_207; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 47:19]
  wire  flags_zf_21 = result_5 == 16'h0; // @[src/main/scala/cpu8086/CPU8086.scala 76:21]
  wire  flags_sf_21 = result_5[15]; // @[src/main/scala/cpu8086/CPU8086.scala 77:20]
  wire [1:0] _flags_pf_T_513 = result_5[0] + result_5[1]; // @[src/main/scala/cpu8086/CPU8086.scala 78:22]
  wire [1:0] _flags_pf_T_515 = result_5[2] + result_5[3]; // @[src/main/scala/cpu8086/CPU8086.scala 78:22]
  wire [2:0] _flags_pf_T_517 = _flags_pf_T_513 + _flags_pf_T_515; // @[src/main/scala/cpu8086/CPU8086.scala 78:22]
  wire [1:0] _flags_pf_T_519 = result_5[4] + result_5[5]; // @[src/main/scala/cpu8086/CPU8086.scala 78:22]
  wire [1:0] _flags_pf_T_521 = result_5[6] + result_5[7]; // @[src/main/scala/cpu8086/CPU8086.scala 78:22]
  wire [2:0] _flags_pf_T_523 = _flags_pf_T_519 + _flags_pf_T_521; // @[src/main/scala/cpu8086/CPU8086.scala 78:22]
  wire [3:0] _flags_pf_T_525 = _flags_pf_T_517 + _flags_pf_T_523; // @[src/main/scala/cpu8086/CPU8086.scala 78:22]
  wire [3:0] _GEN_398 = _flags_pf_T_525 % 4'h2; // @[src/main/scala/cpu8086/CPU8086.scala 78:37]
  wire  flags_pf_21 = _GEN_398[1:0] == 2'h0; // @[src/main/scala/cpu8086/CPU8086.scala 78:43]
  wire [16:0] _flags_T_72 = {9'h0,flags_sf_21,flags_zf_21,1'h0,2'h0,flags_pf_21,2'h0}; // @[src/main/scala/cpu8086/CPU8086.scala 80:8]
  wire [15:0] result_6 = ~srcVal; // @[src/main/scala/cpu8086/CPU8086.scala 300:24]
  wire [15:0] _GEN_216 = _srcVal_T_12 ? result_6 : di; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 118:20 47:19]
  wire [15:0] _GEN_217 = _srcVal_T_10 ? result_6 : si; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 117:20 46:19]
  wire [15:0] _GEN_218 = _srcVal_T_10 ? di : _GEN_216; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 47:19]
  wire [15:0] _GEN_219 = _srcVal_T_8 ? result_6 : bp; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 116:20 45:19]
  wire [15:0] _GEN_220 = _srcVal_T_8 ? si : _GEN_217; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 46:19]
  wire [15:0] _GEN_221 = _srcVal_T_8 ? di : _GEN_218; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 47:19]
  wire [15:0] _GEN_222 = _srcVal_T_6 ? result_6 : sp; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 115:20 44:19]
  wire [15:0] _GEN_223 = _srcVal_T_6 ? bp : _GEN_219; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 45:19]
  wire [15:0] _GEN_224 = _srcVal_T_6 ? si : _GEN_220; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 46:19]
  wire [15:0] _GEN_225 = _srcVal_T_6 ? di : _GEN_221; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 47:19]
  wire [15:0] _GEN_226 = _srcVal_T_4 ? result_6 : bx; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 114:20 41:19]
  wire [15:0] _GEN_227 = _srcVal_T_4 ? sp : _GEN_222; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 44:19]
  wire [15:0] _GEN_228 = _srcVal_T_4 ? bp : _GEN_223; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 45:19]
  wire [15:0] _GEN_229 = _srcVal_T_4 ? si : _GEN_224; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 46:19]
  wire [15:0] _GEN_230 = _srcVal_T_4 ? di : _GEN_225; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 47:19]
  wire [15:0] _GEN_231 = _srcVal_T_2 ? result_6 : dx; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 113:20 43:19]
  wire [15:0] _GEN_232 = _srcVal_T_2 ? bx : _GEN_226; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 41:19]
  wire [15:0] _GEN_233 = _srcVal_T_2 ? sp : _GEN_227; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 44:19]
  wire [15:0] _GEN_234 = _srcVal_T_2 ? bp : _GEN_228; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 45:19]
  wire [15:0] _GEN_235 = _srcVal_T_2 ? si : _GEN_229; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 46:19]
  wire [15:0] _GEN_236 = _srcVal_T_2 ? di : _GEN_230; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 47:19]
  wire [15:0] _GEN_237 = _srcVal_T ? result_6 : cx; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 112:20 42:19]
  wire [15:0] _GEN_238 = _srcVal_T ? dx : _GEN_231; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 43:19]
  wire [15:0] _GEN_239 = _srcVal_T ? bx : _GEN_232; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 41:19]
  wire [15:0] _GEN_240 = _srcVal_T ? sp : _GEN_233; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 44:19]
  wire [15:0] _GEN_241 = _srcVal_T ? bp : _GEN_234; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 45:19]
  wire [15:0] _GEN_242 = _srcVal_T ? si : _GEN_235; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 46:19]
  wire [15:0] _GEN_243 = _srcVal_T ? di : _GEN_236; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 47:19]
  wire [15:0] _GEN_244 = 3'h0 == srcReg ? result_6 : ax; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 111:20 40:19]
  wire [15:0] _GEN_245 = 3'h0 == srcReg ? cx : _GEN_237; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 42:19]
  wire [15:0] _GEN_246 = 3'h0 == srcReg ? dx : _GEN_238; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 43:19]
  wire [15:0] _GEN_247 = 3'h0 == srcReg ? bx : _GEN_239; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 41:19]
  wire [15:0] _GEN_248 = 3'h0 == srcReg ? sp : _GEN_240; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 44:19]
  wire [15:0] _GEN_249 = 3'h0 == srcReg ? bp : _GEN_241; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 45:19]
  wire [15:0] _GEN_250 = 3'h0 == srcReg ? si : _GEN_242; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 46:19]
  wire [15:0] _GEN_251 = 3'h0 == srcReg ? di : _GEN_243; // @[src/main/scala/cpu8086/CPU8086.scala 110:21 47:19]
  wire [15:0] _sp_T_5 = sp - 16'h2; // @[src/main/scala/cpu8086/CPU8086.scala 320:20]
  wire  _T_93 = 8'h58 == opcode; // @[src/main/scala/cpu8086/CPU8086.scala 167:22]
  wire  _T_94 = 8'h59 == opcode; // @[src/main/scala/cpu8086/CPU8086.scala 167:22]
  wire  _T_95 = 8'h5a == opcode; // @[src/main/scala/cpu8086/CPU8086.scala 167:22]
  wire  _T_96 = 8'h5b == opcode; // @[src/main/scala/cpu8086/CPU8086.scala 167:22]
  wire [7:0] _offset_T_2 = operand[7] ? 8'hff : 8'h0; // @[src/main/scala/cpu8086/CPU8086.scala 370:32]
  wire [15:0] offset = {_offset_T_2,operand}; // @[src/main/scala/cpu8086/CPU8086.scala 370:58]
  wire [15:0] _ip_T_6 = $signed(ip) + $signed(offset); // @[src/main/scala/cpu8086/CPU8086.scala 371:38]
  wire  _T_102 = ~flags[6]; // @[src/main/scala/cpu8086/CPU8086.scala 126:23]
  wire  _T_107 = flags[7] == flags[11]; // @[src/main/scala/cpu8086/CPU8086.scala 127:44]
  wire  _T_108 = _T_102 & flags[7] == flags[11]; // @[src/main/scala/cpu8086/CPU8086.scala 127:35]
  wire  _T_111 = flags[7] != flags[11]; // @[src/main/scala/cpu8086/CPU8086.scala 128:23]
  wire  _T_120 = flags[6] | _T_111; // @[src/main/scala/cpu8086/CPU8086.scala 130:34]
  wire [15:0] _GEN_252 = flags[6] ? _ip_T_6 : ip; // @[src/main/scala/cpu8086/CPU8086.scala 377:39 379:16 56:19]
  wire [15:0] _GEN_253 = _T_102 ? _ip_T_6 : ip; // @[src/main/scala/cpu8086/CPU8086.scala 385:39 387:16 56:19]
  wire [15:0] _GEN_254 = _T_108 ? _ip_T_6 : ip; // @[src/main/scala/cpu8086/CPU8086.scala 393:39 395:16 56:19]
  wire [15:0] _GEN_255 = _T_111 ? _ip_T_6 : ip; // @[src/main/scala/cpu8086/CPU8086.scala 401:39 403:16 56:19]
  wire [15:0] _GEN_256 = _T_107 ? _ip_T_6 : ip; // @[src/main/scala/cpu8086/CPU8086.scala 409:39 411:16 56:19]
  wire [15:0] _GEN_257 = _T_120 ? _ip_T_6 : ip; // @[src/main/scala/cpu8086/CPU8086.scala 417:39 419:16 56:19]
  wire  _T_441 = 8'hc3 == opcode; // @[src/main/scala/cpu8086/CPU8086.scala 167:22]
  wire [2:0] _GEN_258 = 8'hf4 == opcode ? 3'h6 : state; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 448:17 61:22]
  wire [2:0] _GEN_259 = 8'h90 == opcode ? 3'h0 : _GEN_258; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 443:17]
  wire [2:0] _GEN_260 = 8'hc3 == opcode ? 3'h5 : _GEN_259; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 436:17]
  wire [15:0] _GEN_262 = 8'he8 == opcode ? _sp_T_5 : sp; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 427:14 44:19]
  wire [15:0] _GEN_263 = 8'he8 == opcode ? ip : memData; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 428:19 64:24]
  wire [15:0] _GEN_264 = 8'he8 == opcode ? _ip_T_6 : ip; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 430:14 56:19]
  wire [2:0] _GEN_265 = 8'he8 == opcode ? 3'h4 : _GEN_260; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 431:17]
  wire [15:0] _GEN_266 = 8'h7e == opcode ? _GEN_257 : _GEN_264; // @[src/main/scala/cpu8086/CPU8086.scala 167:22]
  wire [2:0] _GEN_267 = 8'h7e == opcode ? 3'h0 : _GEN_265; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 421:17]
  wire [15:0] _GEN_269 = 8'h7e == opcode ? sp : _GEN_262; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 44:19]
  wire [15:0] _GEN_270 = 8'h7e == opcode ? memData : _GEN_263; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 64:24]
  wire [15:0] _GEN_271 = 8'h7d == opcode ? _GEN_256 : _GEN_266; // @[src/main/scala/cpu8086/CPU8086.scala 167:22]
  wire [2:0] _GEN_272 = 8'h7d == opcode ? 3'h0 : _GEN_267; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 413:17]
  wire [15:0] _GEN_274 = 8'h7d == opcode ? sp : _GEN_269; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 44:19]
  wire [15:0] _GEN_275 = 8'h7d == opcode ? memData : _GEN_270; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 64:24]
  wire [15:0] _GEN_276 = 8'h7c == opcode ? _GEN_255 : _GEN_271; // @[src/main/scala/cpu8086/CPU8086.scala 167:22]
  wire [2:0] _GEN_277 = 8'h7c == opcode ? 3'h0 : _GEN_272; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 405:17]
  wire [15:0] _GEN_279 = 8'h7c == opcode ? sp : _GEN_274; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 44:19]
  wire [15:0] _GEN_280 = 8'h7c == opcode ? memData : _GEN_275; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 64:24]
  wire [15:0] _GEN_281 = 8'h7f == opcode ? _GEN_254 : _GEN_276; // @[src/main/scala/cpu8086/CPU8086.scala 167:22]
  wire [2:0] _GEN_282 = 8'h7f == opcode ? 3'h0 : _GEN_277; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 397:17]
  wire [15:0] _GEN_284 = 8'h7f == opcode ? sp : _GEN_279; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 44:19]
  wire [15:0] _GEN_285 = 8'h7f == opcode ? memData : _GEN_280; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 64:24]
  wire [15:0] _GEN_286 = 8'h75 == opcode ? _GEN_253 : _GEN_281; // @[src/main/scala/cpu8086/CPU8086.scala 167:22]
  wire [2:0] _GEN_287 = 8'h75 == opcode ? 3'h0 : _GEN_282; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 389:17]
  wire [15:0] _GEN_289 = 8'h75 == opcode ? sp : _GEN_284; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 44:19]
  wire [15:0] _GEN_290 = 8'h75 == opcode ? memData : _GEN_285; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 64:24]
  wire [15:0] _GEN_291 = 8'h74 == opcode ? _GEN_252 : _GEN_286; // @[src/main/scala/cpu8086/CPU8086.scala 167:22]
  wire [2:0] _GEN_292 = 8'h74 == opcode ? 3'h0 : _GEN_287; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 381:17]
  wire [15:0] _GEN_294 = 8'h74 == opcode ? sp : _GEN_289; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 44:19]
  wire [15:0] _GEN_295 = 8'h74 == opcode ? memData : _GEN_290; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 64:24]
  wire [15:0] _GEN_296 = 8'heb == opcode ? _ip_T_6 : _GEN_291; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 371:14]
  wire [2:0] _GEN_297 = 8'heb == opcode ? 3'h0 : _GEN_292; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 372:17]
  wire [15:0] _GEN_299 = 8'heb == opcode ? sp : _GEN_294; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 44:19]
  wire [15:0] _GEN_300 = 8'heb == opcode ? memData : _GEN_295; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 64:24]
  wire [2:0] _GEN_301 = 8'h5b == opcode ? 3'h5 : _GEN_297; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 363:17]
  wire [15:0] _GEN_302 = 8'h5b == opcode ? ip : _GEN_296; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 56:19]
  wire [15:0] _GEN_304 = 8'h5b == opcode ? sp : _GEN_299; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 44:19]
  wire [15:0] _GEN_305 = 8'h5b == opcode ? memData : _GEN_300; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 64:24]
  wire [2:0] _GEN_306 = 8'h5a == opcode ? 3'h5 : _GEN_301; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 358:17]
  wire [15:0] _GEN_307 = 8'h5a == opcode ? ip : _GEN_302; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 56:19]
  wire [15:0] _GEN_309 = 8'h5a == opcode ? sp : _GEN_304; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 44:19]
  wire [15:0] _GEN_310 = 8'h5a == opcode ? memData : _GEN_305; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 64:24]
  wire [2:0] _GEN_311 = 8'h59 == opcode ? 3'h5 : _GEN_306; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 353:17]
  wire [15:0] _GEN_312 = 8'h59 == opcode ? ip : _GEN_307; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 56:19]
  wire [15:0] _GEN_314 = 8'h59 == opcode ? sp : _GEN_309; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 44:19]
  wire [15:0] _GEN_315 = 8'h59 == opcode ? memData : _GEN_310; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 64:24]
  wire [2:0] _GEN_316 = 8'h58 == opcode ? 3'h5 : _GEN_311; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 348:17]
  wire [15:0] _GEN_317 = 8'h58 == opcode ? ip : _GEN_312; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 56:19]
  wire [15:0] _GEN_319 = 8'h58 == opcode ? sp : _GEN_314; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 44:19]
  wire [15:0] _GEN_320 = 8'h58 == opcode ? memData : _GEN_315; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 64:24]
  wire [15:0] _GEN_321 = 8'h53 == opcode ? _sp_T_5 : _GEN_319; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 341:14]
  wire [15:0] _GEN_322 = 8'h53 == opcode ? bx : _GEN_320; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 342:19]
  wire [2:0] _GEN_323 = 8'h53 == opcode ? 3'h4 : _GEN_316; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 343:17]
  wire [15:0] _GEN_324 = 8'h53 == opcode ? ip : _GEN_317; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 56:19]
  wire [15:0] _GEN_326 = 8'h52 == opcode ? _sp_T_5 : _GEN_321; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 334:14]
  wire [15:0] _GEN_327 = 8'h52 == opcode ? dx : _GEN_322; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 335:19]
  wire [2:0] _GEN_328 = 8'h52 == opcode ? 3'h4 : _GEN_323; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 336:17]
  wire [15:0] _GEN_329 = 8'h52 == opcode ? ip : _GEN_324; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 56:19]
  wire [15:0] _GEN_331 = 8'h51 == opcode ? _sp_T_5 : _GEN_326; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 327:14]
  wire [15:0] _GEN_332 = 8'h51 == opcode ? cx : _GEN_327; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 328:19]
  wire [2:0] _GEN_333 = 8'h51 == opcode ? 3'h4 : _GEN_328; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 329:17]
  wire [15:0] _GEN_334 = 8'h51 == opcode ? ip : _GEN_329; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 56:19]
  wire [15:0] _GEN_336 = 8'h50 == opcode ? _sp_T_5 : _GEN_331; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 320:14]
  wire [15:0] _GEN_337 = 8'h50 == opcode ? ax : _GEN_332; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 321:19]
  wire [2:0] _GEN_338 = 8'h50 == opcode ? 3'h4 : _GEN_333; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 322:17]
  wire [15:0] _GEN_339 = 8'h50 == opcode ? ip : _GEN_334; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 56:19]
  wire [16:0] _GEN_341 = 8'h85 == opcode ? _flags_T_70 : {{1'd0}, flags}; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 312:17 57:22]
  wire [2:0] _GEN_342 = 8'h85 == opcode ? 3'h0 : _GEN_338; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 313:17]
  wire [15:0] _GEN_343 = 8'h85 == opcode ? sp : _GEN_336; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 44:19]
  wire [15:0] _GEN_344 = 8'h85 == opcode ? memData : _GEN_337; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 64:24]
  wire [15:0] _GEN_345 = 8'h85 == opcode ? ip : _GEN_339; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 56:19]
  wire [15:0] _GEN_347 = 8'hf7 == opcode ? _GEN_244 : ax; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 40:19]
  wire [15:0] _GEN_348 = 8'hf7 == opcode ? _GEN_245 : cx; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 42:19]
  wire [15:0] _GEN_349 = 8'hf7 == opcode ? _GEN_246 : dx; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 43:19]
  wire [15:0] _GEN_350 = 8'hf7 == opcode ? _GEN_247 : bx; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 41:19]
  wire [15:0] _GEN_351 = 8'hf7 == opcode ? _GEN_248 : _GEN_343; // @[src/main/scala/cpu8086/CPU8086.scala 167:22]
  wire [15:0] _GEN_352 = 8'hf7 == opcode ? _GEN_249 : bp; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 45:19]
  wire [15:0] _GEN_353 = 8'hf7 == opcode ? _GEN_250 : si; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 46:19]
  wire [15:0] _GEN_354 = 8'hf7 == opcode ? _GEN_251 : di; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 47:19]
  wire [2:0] _GEN_355 = 8'hf7 == opcode ? 3'h0 : _GEN_342; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 303:17]
  wire [16:0] _GEN_356 = 8'hf7 == opcode ? {{1'd0}, flags} : _GEN_341; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 57:22]
  wire [15:0] _GEN_357 = 8'hf7 == opcode ? memData : _GEN_344; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 64:24]
  wire [15:0] _GEN_358 = 8'hf7 == opcode ? ip : _GEN_345; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 56:19]
  wire [15:0] _GEN_360 = 8'h31 == opcode ? _GEN_208 : _GEN_347; // @[src/main/scala/cpu8086/CPU8086.scala 167:22]
  wire [15:0] _GEN_361 = 8'h31 == opcode ? _GEN_209 : _GEN_348; // @[src/main/scala/cpu8086/CPU8086.scala 167:22]
  wire [15:0] _GEN_362 = 8'h31 == opcode ? _GEN_210 : _GEN_349; // @[src/main/scala/cpu8086/CPU8086.scala 167:22]
  wire [15:0] _GEN_363 = 8'h31 == opcode ? _GEN_211 : _GEN_350; // @[src/main/scala/cpu8086/CPU8086.scala 167:22]
  wire [15:0] _GEN_364 = 8'h31 == opcode ? _GEN_212 : _GEN_351; // @[src/main/scala/cpu8086/CPU8086.scala 167:22]
  wire [15:0] _GEN_365 = 8'h31 == opcode ? _GEN_213 : _GEN_352; // @[src/main/scala/cpu8086/CPU8086.scala 167:22]
  wire [15:0] _GEN_366 = 8'h31 == opcode ? _GEN_214 : _GEN_353; // @[src/main/scala/cpu8086/CPU8086.scala 167:22]
  wire [15:0] _GEN_367 = 8'h31 == opcode ? _GEN_215 : _GEN_354; // @[src/main/scala/cpu8086/CPU8086.scala 167:22]
  wire [16:0] _GEN_368 = 8'h31 == opcode ? _flags_T_72 : _GEN_356; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 292:17]
  wire [2:0] _GEN_369 = 8'h31 == opcode ? 3'h0 : _GEN_355; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 293:17]
  wire [15:0] _GEN_370 = 8'h31 == opcode ? memData : _GEN_357; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 64:24]
  wire [15:0] _GEN_371 = 8'h31 == opcode ? ip : _GEN_358; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 56:19]
  wire [15:0] _GEN_373 = 8'h9 == opcode ? _GEN_172 : _GEN_360; // @[src/main/scala/cpu8086/CPU8086.scala 167:22]
  wire [15:0] _GEN_374 = 8'h9 == opcode ? _GEN_173 : _GEN_361; // @[src/main/scala/cpu8086/CPU8086.scala 167:22]
  wire [15:0] _GEN_375 = 8'h9 == opcode ? _GEN_174 : _GEN_362; // @[src/main/scala/cpu8086/CPU8086.scala 167:22]
  wire [15:0] _GEN_376 = 8'h9 == opcode ? _GEN_175 : _GEN_363; // @[src/main/scala/cpu8086/CPU8086.scala 167:22]
  wire [15:0] _GEN_377 = 8'h9 == opcode ? _GEN_176 : _GEN_364; // @[src/main/scala/cpu8086/CPU8086.scala 167:22]
  wire [15:0] _GEN_378 = 8'h9 == opcode ? _GEN_177 : _GEN_365; // @[src/main/scala/cpu8086/CPU8086.scala 167:22]
  wire [15:0] _GEN_379 = 8'h9 == opcode ? _GEN_178 : _GEN_366; // @[src/main/scala/cpu8086/CPU8086.scala 167:22]
  wire [15:0] _GEN_380 = 8'h9 == opcode ? _GEN_179 : _GEN_367; // @[src/main/scala/cpu8086/CPU8086.scala 167:22]
  wire [16:0] _GEN_381 = 8'h9 == opcode ? _flags_T_71 : _GEN_368; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 281:17]
  wire [2:0] _GEN_382 = 8'h9 == opcode ? 3'h0 : _GEN_369; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 282:17]
  wire [15:0] _GEN_383 = 8'h9 == opcode ? memData : _GEN_370; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 64:24]
  wire [15:0] _GEN_384 = 8'h9 == opcode ? ip : _GEN_371; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 56:19]
  wire [15:0] _GEN_386 = 8'h21 == opcode ? _GEN_136 : _GEN_373; // @[src/main/scala/cpu8086/CPU8086.scala 167:22]
  wire [15:0] _GEN_387 = 8'h21 == opcode ? _GEN_137 : _GEN_374; // @[src/main/scala/cpu8086/CPU8086.scala 167:22]
  wire [15:0] _GEN_388 = 8'h21 == opcode ? _GEN_138 : _GEN_375; // @[src/main/scala/cpu8086/CPU8086.scala 167:22]
  wire [15:0] _GEN_389 = 8'h21 == opcode ? _GEN_139 : _GEN_376; // @[src/main/scala/cpu8086/CPU8086.scala 167:22]
  wire [15:0] _GEN_390 = 8'h21 == opcode ? _GEN_140 : _GEN_377; // @[src/main/scala/cpu8086/CPU8086.scala 167:22]
  wire [15:0] _GEN_391 = 8'h21 == opcode ? _GEN_141 : _GEN_378; // @[src/main/scala/cpu8086/CPU8086.scala 167:22]
  wire [15:0] _GEN_392 = 8'h21 == opcode ? _GEN_142 : _GEN_379; // @[src/main/scala/cpu8086/CPU8086.scala 167:22]
  wire [15:0] _GEN_393 = 8'h21 == opcode ? _GEN_143 : _GEN_380; // @[src/main/scala/cpu8086/CPU8086.scala 167:22]
  wire [16:0] _GEN_394 = 8'h21 == opcode ? _flags_T_70 : _GEN_381; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 270:17]
  wire [2:0] _GEN_395 = 8'h21 == opcode ? 3'h0 : _GEN_382; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 271:17]
  wire [15:0] _GEN_396 = 8'h21 == opcode ? memData : _GEN_383; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 64:24]
  wire [15:0] _GEN_397 = 8'h21 == opcode ? ip : _GEN_384; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 56:19]
  wire [16:0] _GEN_399 = 8'h39 == opcode ? _flags_T_3 : _GEN_394; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 257:17]
  wire [2:0] _GEN_400 = 8'h39 == opcode ? 3'h0 : _GEN_395; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 258:17]
  wire [15:0] _GEN_401 = 8'h39 == opcode ? ax : _GEN_386; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 40:19]
  wire [15:0] _GEN_402 = 8'h39 == opcode ? cx : _GEN_387; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 42:19]
  wire [15:0] _GEN_403 = 8'h39 == opcode ? dx : _GEN_388; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 43:19]
  wire [15:0] _GEN_404 = 8'h39 == opcode ? bx : _GEN_389; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 41:19]
  wire [15:0] _GEN_405 = 8'h39 == opcode ? sp : _GEN_390; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 44:19]
  wire [15:0] _GEN_406 = 8'h39 == opcode ? bp : _GEN_391; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 45:19]
  wire [15:0] _GEN_407 = 8'h39 == opcode ? si : _GEN_392; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 46:19]
  wire [15:0] _GEN_408 = 8'h39 == opcode ? di : _GEN_393; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 47:19]
  wire [15:0] _GEN_409 = 8'h39 == opcode ? memData : _GEN_396; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 64:24]
  wire [15:0] _GEN_410 = 8'h39 == opcode ? ip : _GEN_397; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 56:19]
  wire [15:0] _GEN_412 = 8'h4f == opcode ? _di_T_3 : _GEN_408; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 247:25]
  wire [16:0] _GEN_413 = 8'h4f == opcode ? _flags_T_67 : _GEN_399; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 247:44]
  wire [2:0] _GEN_414 = 8'h4f == opcode ? 3'h0 : _GEN_400; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 247:92]
  wire [15:0] _GEN_415 = 8'h4f == opcode ? ax : _GEN_401; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 40:19]
  wire [15:0] _GEN_416 = 8'h4f == opcode ? cx : _GEN_402; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 42:19]
  wire [15:0] _GEN_417 = 8'h4f == opcode ? dx : _GEN_403; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 43:19]
  wire [15:0] _GEN_418 = 8'h4f == opcode ? bx : _GEN_404; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 41:19]
  wire [15:0] _GEN_419 = 8'h4f == opcode ? sp : _GEN_405; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 44:19]
  wire [15:0] _GEN_420 = 8'h4f == opcode ? bp : _GEN_406; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 45:19]
  wire [15:0] _GEN_421 = 8'h4f == opcode ? si : _GEN_407; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 46:19]
  wire [15:0] _GEN_422 = 8'h4f == opcode ? memData : _GEN_409; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 64:24]
  wire [15:0] _GEN_423 = 8'h4f == opcode ? ip : _GEN_410; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 56:19]
  wire [15:0] _GEN_425 = 8'h4e == opcode ? _si_T_3 : _GEN_421; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 246:25]
  wire [16:0] _GEN_426 = 8'h4e == opcode ? _flags_T_63 : _GEN_413; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 246:44]
  wire [2:0] _GEN_427 = 8'h4e == opcode ? 3'h0 : _GEN_414; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 246:92]
  wire [15:0] _GEN_428 = 8'h4e == opcode ? di : _GEN_412; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 47:19]
  wire [15:0] _GEN_429 = 8'h4e == opcode ? ax : _GEN_415; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 40:19]
  wire [15:0] _GEN_430 = 8'h4e == opcode ? cx : _GEN_416; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 42:19]
  wire [15:0] _GEN_431 = 8'h4e == opcode ? dx : _GEN_417; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 43:19]
  wire [15:0] _GEN_432 = 8'h4e == opcode ? bx : _GEN_418; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 41:19]
  wire [15:0] _GEN_433 = 8'h4e == opcode ? sp : _GEN_419; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 44:19]
  wire [15:0] _GEN_434 = 8'h4e == opcode ? bp : _GEN_420; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 45:19]
  wire [15:0] _GEN_435 = 8'h4e == opcode ? memData : _GEN_422; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 64:24]
  wire [15:0] _GEN_436 = 8'h4e == opcode ? ip : _GEN_423; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 56:19]
  wire [15:0] _GEN_438 = 8'h4d == opcode ? _bp_T_3 : _GEN_434; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 245:25]
  wire [16:0] _GEN_439 = 8'h4d == opcode ? _flags_T_59 : _GEN_426; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 245:44]
  wire [2:0] _GEN_440 = 8'h4d == opcode ? 3'h0 : _GEN_427; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 245:92]
  wire [15:0] _GEN_441 = 8'h4d == opcode ? si : _GEN_425; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 46:19]
  wire [15:0] _GEN_442 = 8'h4d == opcode ? di : _GEN_428; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 47:19]
  wire [15:0] _GEN_443 = 8'h4d == opcode ? ax : _GEN_429; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 40:19]
  wire [15:0] _GEN_444 = 8'h4d == opcode ? cx : _GEN_430; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 42:19]
  wire [15:0] _GEN_445 = 8'h4d == opcode ? dx : _GEN_431; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 43:19]
  wire [15:0] _GEN_446 = 8'h4d == opcode ? bx : _GEN_432; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 41:19]
  wire [15:0] _GEN_447 = 8'h4d == opcode ? sp : _GEN_433; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 44:19]
  wire [15:0] _GEN_448 = 8'h4d == opcode ? memData : _GEN_435; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 64:24]
  wire [15:0] _GEN_449 = 8'h4d == opcode ? ip : _GEN_436; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 56:19]
  wire [15:0] _GEN_451 = 8'h4c == opcode ? _sp_T_3 : _GEN_447; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 244:25]
  wire [16:0] _GEN_452 = 8'h4c == opcode ? _flags_T_55 : _GEN_439; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 244:44]
  wire [2:0] _GEN_453 = 8'h4c == opcode ? 3'h0 : _GEN_440; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 244:92]
  wire [15:0] _GEN_454 = 8'h4c == opcode ? bp : _GEN_438; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 45:19]
  wire [15:0] _GEN_455 = 8'h4c == opcode ? si : _GEN_441; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 46:19]
  wire [15:0] _GEN_456 = 8'h4c == opcode ? di : _GEN_442; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 47:19]
  wire [15:0] _GEN_457 = 8'h4c == opcode ? ax : _GEN_443; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 40:19]
  wire [15:0] _GEN_458 = 8'h4c == opcode ? cx : _GEN_444; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 42:19]
  wire [15:0] _GEN_459 = 8'h4c == opcode ? dx : _GEN_445; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 43:19]
  wire [15:0] _GEN_460 = 8'h4c == opcode ? bx : _GEN_446; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 41:19]
  wire [15:0] _GEN_461 = 8'h4c == opcode ? memData : _GEN_448; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 64:24]
  wire [15:0] _GEN_462 = 8'h4c == opcode ? ip : _GEN_449; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 56:19]
  wire [15:0] _GEN_464 = 8'h4b == opcode ? _bx_T_4 : _GEN_460; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 243:25]
  wire [16:0] _GEN_465 = 8'h4b == opcode ? _flags_T_51 : _GEN_452; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 243:44]
  wire [2:0] _GEN_466 = 8'h4b == opcode ? 3'h0 : _GEN_453; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 243:92]
  wire [15:0] _GEN_467 = 8'h4b == opcode ? sp : _GEN_451; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 44:19]
  wire [15:0] _GEN_468 = 8'h4b == opcode ? bp : _GEN_454; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 45:19]
  wire [15:0] _GEN_469 = 8'h4b == opcode ? si : _GEN_455; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 46:19]
  wire [15:0] _GEN_470 = 8'h4b == opcode ? di : _GEN_456; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 47:19]
  wire [15:0] _GEN_471 = 8'h4b == opcode ? ax : _GEN_457; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 40:19]
  wire [15:0] _GEN_472 = 8'h4b == opcode ? cx : _GEN_458; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 42:19]
  wire [15:0] _GEN_473 = 8'h4b == opcode ? dx : _GEN_459; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 43:19]
  wire [15:0] _GEN_474 = 8'h4b == opcode ? memData : _GEN_461; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 64:24]
  wire [15:0] _GEN_475 = 8'h4b == opcode ? ip : _GEN_462; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 56:19]
  wire [15:0] _GEN_477 = 8'h4a == opcode ? _dx_T_4 : _GEN_473; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 242:25]
  wire [16:0] _GEN_478 = 8'h4a == opcode ? _flags_T_47 : _GEN_465; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 242:44]
  wire [2:0] _GEN_479 = 8'h4a == opcode ? 3'h0 : _GEN_466; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 242:92]
  wire [15:0] _GEN_480 = 8'h4a == opcode ? bx : _GEN_464; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 41:19]
  wire [15:0] _GEN_481 = 8'h4a == opcode ? sp : _GEN_467; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 44:19]
  wire [15:0] _GEN_482 = 8'h4a == opcode ? bp : _GEN_468; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 45:19]
  wire [15:0] _GEN_483 = 8'h4a == opcode ? si : _GEN_469; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 46:19]
  wire [15:0] _GEN_484 = 8'h4a == opcode ? di : _GEN_470; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 47:19]
  wire [15:0] _GEN_485 = 8'h4a == opcode ? ax : _GEN_471; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 40:19]
  wire [15:0] _GEN_486 = 8'h4a == opcode ? cx : _GEN_472; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 42:19]
  wire [15:0] _GEN_487 = 8'h4a == opcode ? memData : _GEN_474; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 64:24]
  wire [15:0] _GEN_488 = 8'h4a == opcode ? ip : _GEN_475; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 56:19]
  wire [15:0] _GEN_490 = 8'h49 == opcode ? _cx_T_4 : _GEN_486; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 241:25]
  wire [16:0] _GEN_491 = 8'h49 == opcode ? _flags_T_43 : _GEN_478; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 241:44]
  wire [2:0] _GEN_492 = 8'h49 == opcode ? 3'h0 : _GEN_479; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 241:92]
  wire [15:0] _GEN_493 = 8'h49 == opcode ? dx : _GEN_477; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 43:19]
  wire [15:0] _GEN_494 = 8'h49 == opcode ? bx : _GEN_480; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 41:19]
  wire [15:0] _GEN_495 = 8'h49 == opcode ? sp : _GEN_481; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 44:19]
  wire [15:0] _GEN_496 = 8'h49 == opcode ? bp : _GEN_482; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 45:19]
  wire [15:0] _GEN_497 = 8'h49 == opcode ? si : _GEN_483; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 46:19]
  wire [15:0] _GEN_498 = 8'h49 == opcode ? di : _GEN_484; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 47:19]
  wire [15:0] _GEN_499 = 8'h49 == opcode ? ax : _GEN_485; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 40:19]
  wire [15:0] _GEN_500 = 8'h49 == opcode ? memData : _GEN_487; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 64:24]
  wire [15:0] _GEN_501 = 8'h49 == opcode ? ip : _GEN_488; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 56:19]
  wire [15:0] _GEN_503 = 8'h48 == opcode ? _ax_T_4 : _GEN_499; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 240:25]
  wire [16:0] _GEN_504 = 8'h48 == opcode ? _flags_T_39 : _GEN_491; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 240:44]
  wire [2:0] _GEN_505 = 8'h48 == opcode ? 3'h0 : _GEN_492; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 240:92]
  wire [15:0] _GEN_506 = 8'h48 == opcode ? cx : _GEN_490; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 42:19]
  wire [15:0] _GEN_507 = 8'h48 == opcode ? dx : _GEN_493; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 43:19]
  wire [15:0] _GEN_508 = 8'h48 == opcode ? bx : _GEN_494; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 41:19]
  wire [15:0] _GEN_509 = 8'h48 == opcode ? sp : _GEN_495; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 44:19]
  wire [15:0] _GEN_510 = 8'h48 == opcode ? bp : _GEN_496; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 45:19]
  wire [15:0] _GEN_511 = 8'h48 == opcode ? si : _GEN_497; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 46:19]
  wire [15:0] _GEN_512 = 8'h48 == opcode ? di : _GEN_498; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 47:19]
  wire [15:0] _GEN_513 = 8'h48 == opcode ? memData : _GEN_500; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 64:24]
  wire [15:0] _GEN_514 = 8'h48 == opcode ? ip : _GEN_501; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 56:19]
  wire [15:0] _GEN_516 = 8'h47 == opcode ? _di_T_1 : _GEN_512; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 237:25]
  wire [16:0] _GEN_517 = 8'h47 == opcode ? _flags_T_35 : _GEN_504; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 237:44]
  wire [2:0] _GEN_518 = 8'h47 == opcode ? 3'h0 : _GEN_505; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 237:92]
  wire [15:0] _GEN_519 = 8'h47 == opcode ? ax : _GEN_503; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 40:19]
  wire [15:0] _GEN_520 = 8'h47 == opcode ? cx : _GEN_506; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 42:19]
  wire [15:0] _GEN_521 = 8'h47 == opcode ? dx : _GEN_507; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 43:19]
  wire [15:0] _GEN_522 = 8'h47 == opcode ? bx : _GEN_508; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 41:19]
  wire [15:0] _GEN_523 = 8'h47 == opcode ? sp : _GEN_509; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 44:19]
  wire [15:0] _GEN_524 = 8'h47 == opcode ? bp : _GEN_510; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 45:19]
  wire [15:0] _GEN_525 = 8'h47 == opcode ? si : _GEN_511; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 46:19]
  wire [15:0] _GEN_526 = 8'h47 == opcode ? memData : _GEN_513; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 64:24]
  wire [15:0] _GEN_527 = 8'h47 == opcode ? ip : _GEN_514; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 56:19]
  wire [15:0] _GEN_529 = 8'h46 == opcode ? _si_T_1 : _GEN_525; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 236:25]
  wire [16:0] _GEN_530 = 8'h46 == opcode ? _flags_T_31 : _GEN_517; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 236:44]
  wire [2:0] _GEN_531 = 8'h46 == opcode ? 3'h0 : _GEN_518; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 236:92]
  wire [15:0] _GEN_532 = 8'h46 == opcode ? di : _GEN_516; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 47:19]
  wire [15:0] _GEN_533 = 8'h46 == opcode ? ax : _GEN_519; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 40:19]
  wire [15:0] _GEN_534 = 8'h46 == opcode ? cx : _GEN_520; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 42:19]
  wire [15:0] _GEN_535 = 8'h46 == opcode ? dx : _GEN_521; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 43:19]
  wire [15:0] _GEN_536 = 8'h46 == opcode ? bx : _GEN_522; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 41:19]
  wire [15:0] _GEN_537 = 8'h46 == opcode ? sp : _GEN_523; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 44:19]
  wire [15:0] _GEN_538 = 8'h46 == opcode ? bp : _GEN_524; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 45:19]
  wire [15:0] _GEN_539 = 8'h46 == opcode ? memData : _GEN_526; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 64:24]
  wire [15:0] _GEN_540 = 8'h46 == opcode ? ip : _GEN_527; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 56:19]
  wire [15:0] _GEN_542 = 8'h45 == opcode ? _bp_T_1 : _GEN_538; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 235:25]
  wire [16:0] _GEN_543 = 8'h45 == opcode ? _flags_T_27 : _GEN_530; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 235:44]
  wire [2:0] _GEN_544 = 8'h45 == opcode ? 3'h0 : _GEN_531; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 235:92]
  wire [15:0] _GEN_545 = 8'h45 == opcode ? si : _GEN_529; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 46:19]
  wire [15:0] _GEN_546 = 8'h45 == opcode ? di : _GEN_532; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 47:19]
  wire [15:0] _GEN_547 = 8'h45 == opcode ? ax : _GEN_533; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 40:19]
  wire [15:0] _GEN_548 = 8'h45 == opcode ? cx : _GEN_534; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 42:19]
  wire [15:0] _GEN_549 = 8'h45 == opcode ? dx : _GEN_535; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 43:19]
  wire [15:0] _GEN_550 = 8'h45 == opcode ? bx : _GEN_536; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 41:19]
  wire [15:0] _GEN_551 = 8'h45 == opcode ? sp : _GEN_537; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 44:19]
  wire [15:0] _GEN_552 = 8'h45 == opcode ? memData : _GEN_539; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 64:24]
  wire [15:0] _GEN_553 = 8'h45 == opcode ? ip : _GEN_540; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 56:19]
  wire [15:0] _GEN_555 = 8'h44 == opcode ? _sp_T_1 : _GEN_551; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 234:25]
  wire [16:0] _GEN_556 = 8'h44 == opcode ? _flags_T_23 : _GEN_543; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 234:44]
  wire [2:0] _GEN_557 = 8'h44 == opcode ? 3'h0 : _GEN_544; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 234:92]
  wire [15:0] _GEN_558 = 8'h44 == opcode ? bp : _GEN_542; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 45:19]
  wire [15:0] _GEN_559 = 8'h44 == opcode ? si : _GEN_545; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 46:19]
  wire [15:0] _GEN_560 = 8'h44 == opcode ? di : _GEN_546; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 47:19]
  wire [15:0] _GEN_561 = 8'h44 == opcode ? ax : _GEN_547; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 40:19]
  wire [15:0] _GEN_562 = 8'h44 == opcode ? cx : _GEN_548; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 42:19]
  wire [15:0] _GEN_563 = 8'h44 == opcode ? dx : _GEN_549; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 43:19]
  wire [15:0] _GEN_564 = 8'h44 == opcode ? bx : _GEN_550; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 41:19]
  wire [15:0] _GEN_565 = 8'h44 == opcode ? memData : _GEN_552; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 64:24]
  wire [15:0] _GEN_566 = 8'h44 == opcode ? ip : _GEN_553; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 56:19]
  wire [15:0] _GEN_568 = 8'h43 == opcode ? _bx_T_2 : _GEN_564; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 233:25]
  wire [16:0] _GEN_569 = 8'h43 == opcode ? _flags_T_19 : _GEN_556; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 233:44]
  wire [2:0] _GEN_570 = 8'h43 == opcode ? 3'h0 : _GEN_557; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 233:92]
  wire [15:0] _GEN_571 = 8'h43 == opcode ? sp : _GEN_555; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 44:19]
  wire [15:0] _GEN_572 = 8'h43 == opcode ? bp : _GEN_558; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 45:19]
  wire [15:0] _GEN_573 = 8'h43 == opcode ? si : _GEN_559; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 46:19]
  wire [15:0] _GEN_574 = 8'h43 == opcode ? di : _GEN_560; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 47:19]
  wire [15:0] _GEN_575 = 8'h43 == opcode ? ax : _GEN_561; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 40:19]
  wire [15:0] _GEN_576 = 8'h43 == opcode ? cx : _GEN_562; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 42:19]
  wire [15:0] _GEN_577 = 8'h43 == opcode ? dx : _GEN_563; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 43:19]
  wire [15:0] _GEN_578 = 8'h43 == opcode ? memData : _GEN_565; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 64:24]
  wire [15:0] _GEN_579 = 8'h43 == opcode ? ip : _GEN_566; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 56:19]
  wire [15:0] _GEN_581 = 8'h42 == opcode ? _dx_T_2 : _GEN_577; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 232:25]
  wire [16:0] _GEN_582 = 8'h42 == opcode ? _flags_T_15 : _GEN_569; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 232:44]
  wire [2:0] _GEN_583 = 8'h42 == opcode ? 3'h0 : _GEN_570; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 232:92]
  wire [15:0] _GEN_584 = 8'h42 == opcode ? bx : _GEN_568; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 41:19]
  wire [15:0] _GEN_585 = 8'h42 == opcode ? sp : _GEN_571; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 44:19]
  wire [15:0] _GEN_586 = 8'h42 == opcode ? bp : _GEN_572; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 45:19]
  wire [15:0] _GEN_587 = 8'h42 == opcode ? si : _GEN_573; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 46:19]
  wire [15:0] _GEN_588 = 8'h42 == opcode ? di : _GEN_574; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 47:19]
  wire [15:0] _GEN_589 = 8'h42 == opcode ? ax : _GEN_575; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 40:19]
  wire [15:0] _GEN_590 = 8'h42 == opcode ? cx : _GEN_576; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 42:19]
  wire [15:0] _GEN_591 = 8'h42 == opcode ? memData : _GEN_578; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 64:24]
  wire [15:0] _GEN_592 = 8'h42 == opcode ? ip : _GEN_579; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 56:19]
  wire [15:0] _GEN_594 = 8'h41 == opcode ? _cx_T_2 : _GEN_590; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 231:25]
  wire [16:0] _GEN_595 = 8'h41 == opcode ? _flags_T_11 : _GEN_582; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 231:44]
  wire [2:0] _GEN_596 = 8'h41 == opcode ? 3'h0 : _GEN_583; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 231:92]
  wire [15:0] _GEN_597 = 8'h41 == opcode ? dx : _GEN_581; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 43:19]
  wire [15:0] _GEN_598 = 8'h41 == opcode ? bx : _GEN_584; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 41:19]
  wire [15:0] _GEN_599 = 8'h41 == opcode ? sp : _GEN_585; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 44:19]
  wire [15:0] _GEN_600 = 8'h41 == opcode ? bp : _GEN_586; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 45:19]
  wire [15:0] _GEN_601 = 8'h41 == opcode ? si : _GEN_587; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 46:19]
  wire [15:0] _GEN_602 = 8'h41 == opcode ? di : _GEN_588; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 47:19]
  wire [15:0] _GEN_603 = 8'h41 == opcode ? ax : _GEN_589; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 40:19]
  wire [15:0] _GEN_604 = 8'h41 == opcode ? memData : _GEN_591; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 64:24]
  wire [15:0] _GEN_605 = 8'h41 == opcode ? ip : _GEN_592; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 56:19]
  wire [15:0] _GEN_607 = 8'h40 == opcode ? _ax_T_2 : _GEN_603; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 230:25]
  wire [16:0] _GEN_608 = 8'h40 == opcode ? _flags_T_7 : _GEN_595; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 230:44]
  wire [2:0] _GEN_609 = 8'h40 == opcode ? 3'h0 : _GEN_596; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 230:92]
  wire [15:0] _GEN_610 = 8'h40 == opcode ? cx : _GEN_594; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 42:19]
  wire [15:0] _GEN_611 = 8'h40 == opcode ? dx : _GEN_597; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 43:19]
  wire [15:0] _GEN_612 = 8'h40 == opcode ? bx : _GEN_598; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 41:19]
  wire [15:0] _GEN_613 = 8'h40 == opcode ? sp : _GEN_599; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 44:19]
  wire [15:0] _GEN_614 = 8'h40 == opcode ? bp : _GEN_600; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 45:19]
  wire [15:0] _GEN_615 = 8'h40 == opcode ? si : _GEN_601; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 46:19]
  wire [15:0] _GEN_616 = 8'h40 == opcode ? di : _GEN_602; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 47:19]
  wire [15:0] _GEN_617 = 8'h40 == opcode ? memData : _GEN_604; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 64:24]
  wire [15:0] _GEN_618 = 8'h40 == opcode ? ip : _GEN_605; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 56:19]
  wire [15:0] _GEN_620 = 8'h29 == opcode ? _GEN_100 : _GEN_607; // @[src/main/scala/cpu8086/CPU8086.scala 167:22]
  wire [15:0] _GEN_621 = 8'h29 == opcode ? _GEN_101 : _GEN_610; // @[src/main/scala/cpu8086/CPU8086.scala 167:22]
  wire [15:0] _GEN_622 = 8'h29 == opcode ? _GEN_102 : _GEN_611; // @[src/main/scala/cpu8086/CPU8086.scala 167:22]
  wire [15:0] _GEN_623 = 8'h29 == opcode ? _GEN_103 : _GEN_612; // @[src/main/scala/cpu8086/CPU8086.scala 167:22]
  wire [15:0] _GEN_624 = 8'h29 == opcode ? _GEN_104 : _GEN_613; // @[src/main/scala/cpu8086/CPU8086.scala 167:22]
  wire [15:0] _GEN_625 = 8'h29 == opcode ? _GEN_105 : _GEN_614; // @[src/main/scala/cpu8086/CPU8086.scala 167:22]
  wire [15:0] _GEN_626 = 8'h29 == opcode ? _GEN_106 : _GEN_615; // @[src/main/scala/cpu8086/CPU8086.scala 167:22]
  wire [15:0] _GEN_627 = 8'h29 == opcode ? _GEN_107 : _GEN_616; // @[src/main/scala/cpu8086/CPU8086.scala 167:22]
  wire [16:0] _GEN_628 = 8'h29 == opcode ? _flags_T_3 : _GEN_608; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 225:17]
  wire [2:0] _GEN_629 = 8'h29 == opcode ? 3'h0 : _GEN_609; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 226:17]
  wire [15:0] _GEN_630 = 8'h29 == opcode ? memData : _GEN_617; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 64:24]
  wire [15:0] _GEN_631 = 8'h29 == opcode ? ip : _GEN_618; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 56:19]
  wire [15:0] _GEN_633 = 8'h1 == opcode ? _GEN_64 : _GEN_620; // @[src/main/scala/cpu8086/CPU8086.scala 167:22]
  wire [15:0] _GEN_634 = 8'h1 == opcode ? _GEN_65 : _GEN_621; // @[src/main/scala/cpu8086/CPU8086.scala 167:22]
  wire [15:0] _GEN_635 = 8'h1 == opcode ? _GEN_66 : _GEN_622; // @[src/main/scala/cpu8086/CPU8086.scala 167:22]
  wire [15:0] _GEN_636 = 8'h1 == opcode ? _GEN_67 : _GEN_623; // @[src/main/scala/cpu8086/CPU8086.scala 167:22]
  wire [15:0] _GEN_637 = 8'h1 == opcode ? _GEN_68 : _GEN_624; // @[src/main/scala/cpu8086/CPU8086.scala 167:22]
  wire [15:0] _GEN_638 = 8'h1 == opcode ? _GEN_69 : _GEN_625; // @[src/main/scala/cpu8086/CPU8086.scala 167:22]
  wire [15:0] _GEN_639 = 8'h1 == opcode ? _GEN_70 : _GEN_626; // @[src/main/scala/cpu8086/CPU8086.scala 167:22]
  wire [15:0] _GEN_640 = 8'h1 == opcode ? _GEN_71 : _GEN_627; // @[src/main/scala/cpu8086/CPU8086.scala 167:22]
  wire [16:0] _GEN_641 = 8'h1 == opcode ? _flags_T_1 : _GEN_628; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 212:17]
  wire [2:0] _GEN_642 = 8'h1 == opcode ? 3'h0 : _GEN_629; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 213:17]
  wire [15:0] _GEN_643 = 8'h1 == opcode ? memData : _GEN_630; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 64:24]
  wire [15:0] _GEN_644 = 8'h1 == opcode ? ip : _GEN_631; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 56:19]
  wire [15:0] _GEN_646 = 8'hba == opcode ? _ax_T : _GEN_635; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 197:14]
  wire [2:0] _GEN_647 = 8'hba == opcode ? 3'h0 : _GEN_642; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 198:17]
  wire [15:0] _GEN_648 = 8'hba == opcode ? ax : _GEN_633; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 40:19]
  wire [15:0] _GEN_649 = 8'hba == opcode ? cx : _GEN_634; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 42:19]
  wire [15:0] _GEN_650 = 8'hba == opcode ? bx : _GEN_636; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 41:19]
  wire [15:0] _GEN_651 = 8'hba == opcode ? sp : _GEN_637; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 44:19]
  wire [15:0] _GEN_652 = 8'hba == opcode ? bp : _GEN_638; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 45:19]
  wire [15:0] _GEN_653 = 8'hba == opcode ? si : _GEN_639; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 46:19]
  wire [15:0] _GEN_654 = 8'hba == opcode ? di : _GEN_640; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 47:19]
  wire [16:0] _GEN_655 = 8'hba == opcode ? {{1'd0}, flags} : _GEN_641; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 57:22]
  wire [15:0] _GEN_656 = 8'hba == opcode ? memData : _GEN_643; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 64:24]
  wire [15:0] _GEN_657 = 8'hba == opcode ? ip : _GEN_644; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 56:19]
  wire [15:0] _GEN_659 = 8'hb9 == opcode ? _ax_T : _GEN_649; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 191:14]
  wire [2:0] _GEN_660 = 8'hb9 == opcode ? 3'h0 : _GEN_647; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 192:17]
  wire [15:0] _GEN_661 = 8'hb9 == opcode ? dx : _GEN_646; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 43:19]
  wire [15:0] _GEN_662 = 8'hb9 == opcode ? ax : _GEN_648; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 40:19]
  wire [15:0] _GEN_663 = 8'hb9 == opcode ? bx : _GEN_650; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 41:19]
  wire [15:0] _GEN_664 = 8'hb9 == opcode ? sp : _GEN_651; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 44:19]
  wire [15:0] _GEN_665 = 8'hb9 == opcode ? bp : _GEN_652; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 45:19]
  wire [15:0] _GEN_666 = 8'hb9 == opcode ? si : _GEN_653; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 46:19]
  wire [15:0] _GEN_667 = 8'hb9 == opcode ? di : _GEN_654; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 47:19]
  wire [16:0] _GEN_668 = 8'hb9 == opcode ? {{1'd0}, flags} : _GEN_655; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 57:22]
  wire [15:0] _GEN_669 = 8'hb9 == opcode ? memData : _GEN_656; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 64:24]
  wire [15:0] _GEN_670 = 8'hb9 == opcode ? ip : _GEN_657; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 56:19]
  wire [15:0] _GEN_672 = 8'hbb == opcode ? _ax_T : _GEN_663; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 185:14]
  wire [2:0] _GEN_673 = 8'hbb == opcode ? 3'h0 : _GEN_660; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 186:17]
  wire [15:0] _GEN_674 = 8'hbb == opcode ? cx : _GEN_659; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 42:19]
  wire [15:0] _GEN_675 = 8'hbb == opcode ? dx : _GEN_661; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 43:19]
  wire [15:0] _GEN_676 = 8'hbb == opcode ? ax : _GEN_662; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 40:19]
  wire [15:0] _GEN_677 = 8'hbb == opcode ? sp : _GEN_664; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 44:19]
  wire [15:0] _GEN_678 = 8'hbb == opcode ? bp : _GEN_665; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 45:19]
  wire [15:0] _GEN_679 = 8'hbb == opcode ? si : _GEN_666; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 46:19]
  wire [15:0] _GEN_680 = 8'hbb == opcode ? di : _GEN_667; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 47:19]
  wire [16:0] _GEN_681 = 8'hbb == opcode ? {{1'd0}, flags} : _GEN_668; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 57:22]
  wire [15:0] _GEN_682 = 8'hbb == opcode ? memData : _GEN_669; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 64:24]
  wire [15:0] _GEN_683 = 8'hbb == opcode ? ip : _GEN_670; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 56:19]
  wire [15:0] _GEN_685 = 8'hb8 == opcode ? _ax_T : _GEN_676; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 179:14]
  wire [2:0] _GEN_686 = 8'hb8 == opcode ? 3'h0 : _GEN_673; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 180:17]
  wire [15:0] _GEN_687 = 8'hb8 == opcode ? bx : _GEN_672; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 41:19]
  wire [15:0] _GEN_688 = 8'hb8 == opcode ? cx : _GEN_674; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 42:19]
  wire [15:0] _GEN_689 = 8'hb8 == opcode ? dx : _GEN_675; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 43:19]
  wire [15:0] _GEN_690 = 8'hb8 == opcode ? sp : _GEN_677; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 44:19]
  wire [15:0] _GEN_691 = 8'hb8 == opcode ? bp : _GEN_678; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 45:19]
  wire [15:0] _GEN_692 = 8'hb8 == opcode ? si : _GEN_679; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 46:19]
  wire [15:0] _GEN_693 = 8'hb8 == opcode ? di : _GEN_680; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 47:19]
  wire [16:0] _GEN_694 = 8'hb8 == opcode ? {{1'd0}, flags} : _GEN_681; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 57:22]
  wire [15:0] _GEN_695 = 8'hb8 == opcode ? memData : _GEN_682; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 64:24]
  wire [15:0] _GEN_696 = 8'hb8 == opcode ? ip : _GEN_683; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 56:19]
  wire [2:0] _GEN_706 = 8'h89 == opcode ? 3'h0 : _GEN_686; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 174:17]
  wire [16:0] _GEN_707 = 8'h89 == opcode ? {{1'd0}, flags} : _GEN_694; // @[src/main/scala/cpu8086/CPU8086.scala 167:22 57:22]
  wire [19:0] _GEN_789 = {{4'd0}, sp}; // @[src/main/scala/cpu8086/CPU8086.scala 458:31]
  wire [20:0] _io_memAddr_T_7 = {{1'd0}, _GEN_789}; // @[src/main/scala/cpu8086/CPU8086.scala 458:31]
  wire [15:0] _GEN_712 = _T_441 ? io_memDataIn : ip; // @[src/main/scala/cpu8086/CPU8086.scala 471:26 476:25 56:19]
  wire [15:0] _GEN_713 = _T_96 ? io_memDataIn : bx; // @[src/main/scala/cpu8086/CPU8086.scala 41:19 471:26 475:25]
  wire [15:0] _GEN_714 = _T_96 ? ip : _GEN_712; // @[src/main/scala/cpu8086/CPU8086.scala 471:26 56:19]
  wire [15:0] _GEN_715 = _T_95 ? io_memDataIn : dx; // @[src/main/scala/cpu8086/CPU8086.scala 43:19 471:26 474:25]
  wire [15:0] _GEN_716 = _T_95 ? bx : _GEN_713; // @[src/main/scala/cpu8086/CPU8086.scala 41:19 471:26]
  wire [15:0] _GEN_717 = _T_95 ? ip : _GEN_714; // @[src/main/scala/cpu8086/CPU8086.scala 471:26 56:19]
  wire [15:0] _GEN_718 = _T_94 ? io_memDataIn : cx; // @[src/main/scala/cpu8086/CPU8086.scala 42:19 471:26 473:25]
  wire [15:0] _GEN_719 = _T_94 ? dx : _GEN_715; // @[src/main/scala/cpu8086/CPU8086.scala 43:19 471:26]
  wire [15:0] _GEN_720 = _T_94 ? bx : _GEN_716; // @[src/main/scala/cpu8086/CPU8086.scala 41:19 471:26]
  wire [15:0] _GEN_721 = _T_94 ? ip : _GEN_717; // @[src/main/scala/cpu8086/CPU8086.scala 471:26 56:19]
  wire [15:0] _GEN_722 = _T_93 ? io_memDataIn : ax; // @[src/main/scala/cpu8086/CPU8086.scala 40:19 471:26 472:25]
  wire [15:0] _GEN_723 = _T_93 ? cx : _GEN_718; // @[src/main/scala/cpu8086/CPU8086.scala 42:19 471:26]
  wire [15:0] _GEN_724 = _T_93 ? dx : _GEN_719; // @[src/main/scala/cpu8086/CPU8086.scala 43:19 471:26]
  wire [15:0] _GEN_725 = _T_93 ? bx : _GEN_720; // @[src/main/scala/cpu8086/CPU8086.scala 41:19 471:26]
  wire [15:0] _GEN_726 = _T_93 ? ip : _GEN_721; // @[src/main/scala/cpu8086/CPU8086.scala 471:26 56:19]
  wire [15:0] _sp_T_15 = sp + 16'h2; // @[src/main/scala/cpu8086/CPU8086.scala 479:16]
  wire [19:0] _GEN_728 = 3'h5 == state ? _io_memAddr_T_7[19:0] : _io_memAddr_T_2; // @[src/main/scala/cpu8086/CPU8086.scala 139:14 152:17 465:18]
  wire [15:0] _GEN_730 = 3'h5 == state ? _GEN_722 : ax; // @[src/main/scala/cpu8086/CPU8086.scala 152:17 40:19]
  wire [15:0] _GEN_731 = 3'h5 == state ? _GEN_723 : cx; // @[src/main/scala/cpu8086/CPU8086.scala 152:17 42:19]
  wire [15:0] _GEN_732 = 3'h5 == state ? _GEN_724 : dx; // @[src/main/scala/cpu8086/CPU8086.scala 152:17 43:19]
  wire [15:0] _GEN_733 = 3'h5 == state ? _GEN_725 : bx; // @[src/main/scala/cpu8086/CPU8086.scala 152:17 41:19]
  wire [15:0] _GEN_734 = 3'h5 == state ? _GEN_726 : ip; // @[src/main/scala/cpu8086/CPU8086.scala 152:17 56:19]
  wire [15:0] _GEN_735 = 3'h5 == state ? _sp_T_15 : sp; // @[src/main/scala/cpu8086/CPU8086.scala 152:17 479:10 44:19]
  wire [2:0] _GEN_736 = 3'h5 == state ? 3'h0 : state; // @[src/main/scala/cpu8086/CPU8086.scala 152:17 480:13 61:22]
  wire  _GEN_737 = 3'h5 == state ? 1'h0 : 3'h6 == state; // @[src/main/scala/cpu8086/CPU8086.scala 143:11 152:17]
  wire [19:0] _GEN_738 = 3'h4 == state ? _io_memAddr_T_7[19:0] : _GEN_728; // @[src/main/scala/cpu8086/CPU8086.scala 152:17 458:18]
  wire [15:0] _GEN_739 = 3'h4 == state ? memData : 16'h0; // @[src/main/scala/cpu8086/CPU8086.scala 140:17 152:17 459:21]
  wire  _GEN_742 = 3'h4 == state ? 1'h0 : 3'h5 == state; // @[src/main/scala/cpu8086/CPU8086.scala 142:14 152:17]
  wire  _GEN_749 = 3'h4 == state ? 1'h0 : _GEN_737; // @[src/main/scala/cpu8086/CPU8086.scala 143:11 152:17]
  wire [16:0] _GEN_759 = 3'h1 == state ? _GEN_707 : {{1'd0}, flags}; // @[src/main/scala/cpu8086/CPU8086.scala 152:17 57:22]
  wire [19:0] _GEN_763 = 3'h1 == state ? _io_memAddr_T_2 : _GEN_738; // @[src/main/scala/cpu8086/CPU8086.scala 139:14 152:17]
  wire [15:0] _GEN_764 = 3'h1 == state ? 16'h0 : _GEN_739; // @[src/main/scala/cpu8086/CPU8086.scala 140:17 152:17]
  wire  _GEN_765 = 3'h1 == state ? 1'h0 : 3'h4 == state; // @[src/main/scala/cpu8086/CPU8086.scala 141:15 152:17]
  wire  _GEN_766 = 3'h1 == state ? 1'h0 : _GEN_742; // @[src/main/scala/cpu8086/CPU8086.scala 142:14 152:17]
  wire  _GEN_767 = 3'h1 == state ? 1'h0 : _GEN_749; // @[src/main/scala/cpu8086/CPU8086.scala 143:11 152:17]
  wire [16:0] _GEN_781 = 3'h0 == state ? {{1'd0}, flags} : _GEN_759; // @[src/main/scala/cpu8086/CPU8086.scala 152:17 57:22]
  wire [16:0] _GEN_791 = reset ? 17'h0 : _GEN_781; // @[src/main/scala/cpu8086/CPU8086.scala 57:{22,22}]
  assign io_memAddr = 3'h0 == state ? _io_memAddr_T_2 : _GEN_763; // @[src/main/scala/cpu8086/CPU8086.scala 152:17 154:18]
  assign io_memDataOut = 3'h0 == state ? 16'h0 : _GEN_764; // @[src/main/scala/cpu8086/CPU8086.scala 140:17 152:17]
  assign io_memWrite = 3'h0 == state ? 1'h0 : _GEN_765; // @[src/main/scala/cpu8086/CPU8086.scala 141:15 152:17]
  assign io_memRead = 3'h0 == state | _GEN_766; // @[src/main/scala/cpu8086/CPU8086.scala 152:17 155:18]
  assign io_halt = 3'h0 == state ? 1'h0 : _GEN_767; // @[src/main/scala/cpu8086/CPU8086.scala 143:11 152:17]
  assign io_ax = ax; // @[src/main/scala/cpu8086/CPU8086.scala 144:9]
  assign io_bx = bx; // @[src/main/scala/cpu8086/CPU8086.scala 145:9]
  assign io_cx = cx; // @[src/main/scala/cpu8086/CPU8086.scala 146:9]
  assign io_dx = dx; // @[src/main/scala/cpu8086/CPU8086.scala 147:9]
  assign io_sp = sp; // @[src/main/scala/cpu8086/CPU8086.scala 148:9]
  assign io_ip = ip; // @[src/main/scala/cpu8086/CPU8086.scala 149:9]
  assign io_flags = flags; // @[src/main/scala/cpu8086/CPU8086.scala 150:12]
  always @(posedge clock) begin
    if (reset) begin // @[src/main/scala/cpu8086/CPU8086.scala 40:19]
      ax <= 16'h0; // @[src/main/scala/cpu8086/CPU8086.scala 40:19]
    end else if (!(3'h0 == state)) begin // @[src/main/scala/cpu8086/CPU8086.scala 152:17]
      if (3'h1 == state) begin // @[src/main/scala/cpu8086/CPU8086.scala 152:17]
        if (8'h89 == opcode) begin // @[src/main/scala/cpu8086/CPU8086.scala 167:22]
          ax <= _GEN_28;
        end else begin
          ax <= _GEN_685;
        end
      end else if (!(3'h4 == state)) begin // @[src/main/scala/cpu8086/CPU8086.scala 152:17]
        ax <= _GEN_730;
      end
    end
    if (reset) begin // @[src/main/scala/cpu8086/CPU8086.scala 41:19]
      bx <= 16'h0; // @[src/main/scala/cpu8086/CPU8086.scala 41:19]
    end else if (!(3'h0 == state)) begin // @[src/main/scala/cpu8086/CPU8086.scala 152:17]
      if (3'h1 == state) begin // @[src/main/scala/cpu8086/CPU8086.scala 152:17]
        if (8'h89 == opcode) begin // @[src/main/scala/cpu8086/CPU8086.scala 167:22]
          bx <= _GEN_31;
        end else begin
          bx <= _GEN_687;
        end
      end else if (!(3'h4 == state)) begin // @[src/main/scala/cpu8086/CPU8086.scala 152:17]
        bx <= _GEN_733;
      end
    end
    if (reset) begin // @[src/main/scala/cpu8086/CPU8086.scala 42:19]
      cx <= 16'h0; // @[src/main/scala/cpu8086/CPU8086.scala 42:19]
    end else if (!(3'h0 == state)) begin // @[src/main/scala/cpu8086/CPU8086.scala 152:17]
      if (3'h1 == state) begin // @[src/main/scala/cpu8086/CPU8086.scala 152:17]
        if (8'h89 == opcode) begin // @[src/main/scala/cpu8086/CPU8086.scala 167:22]
          cx <= _GEN_29;
        end else begin
          cx <= _GEN_688;
        end
      end else if (!(3'h4 == state)) begin // @[src/main/scala/cpu8086/CPU8086.scala 152:17]
        cx <= _GEN_731;
      end
    end
    if (reset) begin // @[src/main/scala/cpu8086/CPU8086.scala 43:19]
      dx <= 16'h0; // @[src/main/scala/cpu8086/CPU8086.scala 43:19]
    end else if (!(3'h0 == state)) begin // @[src/main/scala/cpu8086/CPU8086.scala 152:17]
      if (3'h1 == state) begin // @[src/main/scala/cpu8086/CPU8086.scala 152:17]
        if (8'h89 == opcode) begin // @[src/main/scala/cpu8086/CPU8086.scala 167:22]
          dx <= _GEN_30;
        end else begin
          dx <= _GEN_689;
        end
      end else if (!(3'h4 == state)) begin // @[src/main/scala/cpu8086/CPU8086.scala 152:17]
        dx <= _GEN_732;
      end
    end
    if (reset) begin // @[src/main/scala/cpu8086/CPU8086.scala 44:19]
      sp <= 16'hfffe; // @[src/main/scala/cpu8086/CPU8086.scala 44:19]
    end else if (!(3'h0 == state)) begin // @[src/main/scala/cpu8086/CPU8086.scala 152:17]
      if (3'h1 == state) begin // @[src/main/scala/cpu8086/CPU8086.scala 152:17]
        if (8'h89 == opcode) begin // @[src/main/scala/cpu8086/CPU8086.scala 167:22]
          sp <= _GEN_32;
        end else begin
          sp <= _GEN_690;
        end
      end else if (!(3'h4 == state)) begin // @[src/main/scala/cpu8086/CPU8086.scala 152:17]
        sp <= _GEN_735;
      end
    end
    if (reset) begin // @[src/main/scala/cpu8086/CPU8086.scala 45:19]
      bp <= 16'h0; // @[src/main/scala/cpu8086/CPU8086.scala 45:19]
    end else if (!(3'h0 == state)) begin // @[src/main/scala/cpu8086/CPU8086.scala 152:17]
      if (3'h1 == state) begin // @[src/main/scala/cpu8086/CPU8086.scala 152:17]
        if (8'h89 == opcode) begin // @[src/main/scala/cpu8086/CPU8086.scala 167:22]
          bp <= _GEN_33;
        end else begin
          bp <= _GEN_691;
        end
      end
    end
    if (reset) begin // @[src/main/scala/cpu8086/CPU8086.scala 46:19]
      si <= 16'h0; // @[src/main/scala/cpu8086/CPU8086.scala 46:19]
    end else if (!(3'h0 == state)) begin // @[src/main/scala/cpu8086/CPU8086.scala 152:17]
      if (3'h1 == state) begin // @[src/main/scala/cpu8086/CPU8086.scala 152:17]
        if (8'h89 == opcode) begin // @[src/main/scala/cpu8086/CPU8086.scala 167:22]
          si <= _GEN_34;
        end else begin
          si <= _GEN_692;
        end
      end
    end
    if (reset) begin // @[src/main/scala/cpu8086/CPU8086.scala 47:19]
      di <= 16'h0; // @[src/main/scala/cpu8086/CPU8086.scala 47:19]
    end else if (!(3'h0 == state)) begin // @[src/main/scala/cpu8086/CPU8086.scala 152:17]
      if (3'h1 == state) begin // @[src/main/scala/cpu8086/CPU8086.scala 152:17]
        if (8'h89 == opcode) begin // @[src/main/scala/cpu8086/CPU8086.scala 167:22]
          di <= _GEN_35;
        end else begin
          di <= _GEN_693;
        end
      end
    end
    if (reset) begin // @[src/main/scala/cpu8086/CPU8086.scala 56:19]
      ip <= 16'h0; // @[src/main/scala/cpu8086/CPU8086.scala 56:19]
    end else if (3'h0 == state) begin // @[src/main/scala/cpu8086/CPU8086.scala 152:17]
      ip <= _ip_T_1; // @[src/main/scala/cpu8086/CPU8086.scala 157:10]
    end else if (3'h1 == state) begin // @[src/main/scala/cpu8086/CPU8086.scala 152:17]
      if (!(8'h89 == opcode)) begin // @[src/main/scala/cpu8086/CPU8086.scala 167:22]
        ip <= _GEN_696;
      end
    end else if (!(3'h4 == state)) begin // @[src/main/scala/cpu8086/CPU8086.scala 152:17]
      ip <= _GEN_734;
    end
    flags <= _GEN_791[15:0]; // @[src/main/scala/cpu8086/CPU8086.scala 57:{22,22}]
    if (reset) begin // @[src/main/scala/cpu8086/CPU8086.scala 61:22]
      state <= 3'h0; // @[src/main/scala/cpu8086/CPU8086.scala 61:22]
    end else if (3'h0 == state) begin // @[src/main/scala/cpu8086/CPU8086.scala 152:17]
      state <= 3'h1; // @[src/main/scala/cpu8086/CPU8086.scala 158:13]
    end else if (3'h1 == state) begin // @[src/main/scala/cpu8086/CPU8086.scala 152:17]
      if (opcode != 8'hf4 & state == 3'h1) begin // @[src/main/scala/cpu8086/CPU8086.scala 452:53]
        state <= 3'h0; // @[src/main/scala/cpu8086/CPU8086.scala 453:15]
      end else begin
        state <= _GEN_706;
      end
    end else if (3'h4 == state) begin // @[src/main/scala/cpu8086/CPU8086.scala 152:17]
      state <= 3'h0; // @[src/main/scala/cpu8086/CPU8086.scala 461:13]
    end else begin
      state <= _GEN_736;
    end
    if (reset) begin // @[src/main/scala/cpu8086/CPU8086.scala 63:28]
      instruction <= 16'h0; // @[src/main/scala/cpu8086/CPU8086.scala 63:28]
    end else if (3'h0 == state) begin // @[src/main/scala/cpu8086/CPU8086.scala 152:17]
      instruction <= io_memDataIn; // @[src/main/scala/cpu8086/CPU8086.scala 156:19]
    end
    if (reset) begin // @[src/main/scala/cpu8086/CPU8086.scala 64:24]
      memData <= 16'h0; // @[src/main/scala/cpu8086/CPU8086.scala 64:24]
    end else if (!(3'h0 == state)) begin // @[src/main/scala/cpu8086/CPU8086.scala 152:17]
      if (3'h1 == state) begin // @[src/main/scala/cpu8086/CPU8086.scala 152:17]
        if (!(8'h89 == opcode)) begin // @[src/main/scala/cpu8086/CPU8086.scala 167:22]
          memData <= _GEN_695;
        end
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ax = _RAND_0[15:0];
  _RAND_1 = {1{`RANDOM}};
  bx = _RAND_1[15:0];
  _RAND_2 = {1{`RANDOM}};
  cx = _RAND_2[15:0];
  _RAND_3 = {1{`RANDOM}};
  dx = _RAND_3[15:0];
  _RAND_4 = {1{`RANDOM}};
  sp = _RAND_4[15:0];
  _RAND_5 = {1{`RANDOM}};
  bp = _RAND_5[15:0];
  _RAND_6 = {1{`RANDOM}};
  si = _RAND_6[15:0];
  _RAND_7 = {1{`RANDOM}};
  di = _RAND_7[15:0];
  _RAND_8 = {1{`RANDOM}};
  ip = _RAND_8[15:0];
  _RAND_9 = {1{`RANDOM}};
  flags = _RAND_9[15:0];
  _RAND_10 = {1{`RANDOM}};
  state = _RAND_10[2:0];
  _RAND_11 = {1{`RANDOM}};
  instruction = _RAND_11[15:0];
  _RAND_12 = {1{`RANDOM}};
  memData = _RAND_12[15:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Memory(
  input         clock,
  input  [19:0] io_addr, // @[src/main/scala/cpu8086/Memory.scala 13:14]
  input  [15:0] io_dataIn, // @[src/main/scala/cpu8086/Memory.scala 13:14]
  output [15:0] io_dataOut, // @[src/main/scala/cpu8086/Memory.scala 13:14]
  input         io_write, // @[src/main/scala/cpu8086/Memory.scala 13:14]
  input         io_read // @[src/main/scala/cpu8086/Memory.scala 13:14]
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [15:0] mem [0:32767]; // @[src/main/scala/cpu8086/Memory.scala 22:24]
  wire  mem_io_dataOut_MPORT_en; // @[src/main/scala/cpu8086/Memory.scala 22:24]
  wire [14:0] mem_io_dataOut_MPORT_addr; // @[src/main/scala/cpu8086/Memory.scala 22:24]
  wire [15:0] mem_io_dataOut_MPORT_data; // @[src/main/scala/cpu8086/Memory.scala 22:24]
  wire [15:0] mem_MPORT_data; // @[src/main/scala/cpu8086/Memory.scala 22:24]
  wire [14:0] mem_MPORT_addr; // @[src/main/scala/cpu8086/Memory.scala 22:24]
  wire  mem_MPORT_mask; // @[src/main/scala/cpu8086/Memory.scala 22:24]
  wire  mem_MPORT_en; // @[src/main/scala/cpu8086/Memory.scala 22:24]
  reg  mem_io_dataOut_MPORT_en_pipe_0;
  reg [14:0] mem_io_dataOut_MPORT_addr_pipe_0;
  assign mem_io_dataOut_MPORT_en = mem_io_dataOut_MPORT_en_pipe_0;
  assign mem_io_dataOut_MPORT_addr = mem_io_dataOut_MPORT_addr_pipe_0;
  assign mem_io_dataOut_MPORT_data = mem[mem_io_dataOut_MPORT_addr]; // @[src/main/scala/cpu8086/Memory.scala 22:24]
  assign mem_MPORT_data = io_dataIn;
  assign mem_MPORT_addr = io_addr[15:1];
  assign mem_MPORT_mask = 1'h1;
  assign mem_MPORT_en = io_write;
  assign io_dataOut = io_read ? mem_io_dataOut_MPORT_data : 16'h0; // @[src/main/scala/cpu8086/Memory.scala 25:14 28:17 29:16]
  always @(posedge clock) begin
    if (mem_MPORT_en & mem_MPORT_mask) begin
      mem[mem_MPORT_addr] <= mem_MPORT_data; // @[src/main/scala/cpu8086/Memory.scala 22:24]
    end
    mem_io_dataOut_MPORT_en_pipe_0 <= io_read;
    if (io_read) begin
      mem_io_dataOut_MPORT_addr_pipe_0 <= io_addr[15:1];
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 32768; initvar = initvar+1)
    mem[initvar] = _RAND_0[15:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  mem_io_dataOut_MPORT_en_pipe_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  mem_io_dataOut_MPORT_addr_pipe_0 = _RAND_2[14:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module MyCPU8086System(
  input         clock,
  input         reset,
  output        io_halt, // @[src/main/scala/cpu8086/CPU8086.scala 491:14]
  output [15:0] io_ax, // @[src/main/scala/cpu8086/CPU8086.scala 491:14]
  output [15:0] io_bx, // @[src/main/scala/cpu8086/CPU8086.scala 491:14]
  output [15:0] io_cx, // @[src/main/scala/cpu8086/CPU8086.scala 491:14]
  output [15:0] io_dx, // @[src/main/scala/cpu8086/CPU8086.scala 491:14]
  output [15:0] io_sp, // @[src/main/scala/cpu8086/CPU8086.scala 491:14]
  output [15:0] io_ip, // @[src/main/scala/cpu8086/CPU8086.scala 491:14]
  output [15:0] io_flags // @[src/main/scala/cpu8086/CPU8086.scala 491:14]
);
  wire  cpu_clock; // @[src/main/scala/cpu8086/CPU8086.scala 502:19]
  wire  cpu_reset; // @[src/main/scala/cpu8086/CPU8086.scala 502:19]
  wire [19:0] cpu_io_memAddr; // @[src/main/scala/cpu8086/CPU8086.scala 502:19]
  wire [15:0] cpu_io_memDataOut; // @[src/main/scala/cpu8086/CPU8086.scala 502:19]
  wire [15:0] cpu_io_memDataIn; // @[src/main/scala/cpu8086/CPU8086.scala 502:19]
  wire  cpu_io_memWrite; // @[src/main/scala/cpu8086/CPU8086.scala 502:19]
  wire  cpu_io_memRead; // @[src/main/scala/cpu8086/CPU8086.scala 502:19]
  wire  cpu_io_halt; // @[src/main/scala/cpu8086/CPU8086.scala 502:19]
  wire [15:0] cpu_io_ax; // @[src/main/scala/cpu8086/CPU8086.scala 502:19]
  wire [15:0] cpu_io_bx; // @[src/main/scala/cpu8086/CPU8086.scala 502:19]
  wire [15:0] cpu_io_cx; // @[src/main/scala/cpu8086/CPU8086.scala 502:19]
  wire [15:0] cpu_io_dx; // @[src/main/scala/cpu8086/CPU8086.scala 502:19]
  wire [15:0] cpu_io_sp; // @[src/main/scala/cpu8086/CPU8086.scala 502:19]
  wire [15:0] cpu_io_ip; // @[src/main/scala/cpu8086/CPU8086.scala 502:19]
  wire [15:0] cpu_io_flags; // @[src/main/scala/cpu8086/CPU8086.scala 502:19]
  wire  mem_clock; // @[src/main/scala/cpu8086/CPU8086.scala 503:19]
  wire [19:0] mem_io_addr; // @[src/main/scala/cpu8086/CPU8086.scala 503:19]
  wire [15:0] mem_io_dataIn; // @[src/main/scala/cpu8086/CPU8086.scala 503:19]
  wire [15:0] mem_io_dataOut; // @[src/main/scala/cpu8086/CPU8086.scala 503:19]
  wire  mem_io_write; // @[src/main/scala/cpu8086/CPU8086.scala 503:19]
  wire  mem_io_read; // @[src/main/scala/cpu8086/CPU8086.scala 503:19]
  MyCPU8086 cpu ( // @[src/main/scala/cpu8086/CPU8086.scala 502:19]
    .clock(cpu_clock),
    .reset(cpu_reset),
    .io_memAddr(cpu_io_memAddr),
    .io_memDataOut(cpu_io_memDataOut),
    .io_memDataIn(cpu_io_memDataIn),
    .io_memWrite(cpu_io_memWrite),
    .io_memRead(cpu_io_memRead),
    .io_halt(cpu_io_halt),
    .io_ax(cpu_io_ax),
    .io_bx(cpu_io_bx),
    .io_cx(cpu_io_cx),
    .io_dx(cpu_io_dx),
    .io_sp(cpu_io_sp),
    .io_ip(cpu_io_ip),
    .io_flags(cpu_io_flags)
  );
  Memory mem ( // @[src/main/scala/cpu8086/CPU8086.scala 503:19]
    .clock(mem_clock),
    .io_addr(mem_io_addr),
    .io_dataIn(mem_io_dataIn),
    .io_dataOut(mem_io_dataOut),
    .io_write(mem_io_write),
    .io_read(mem_io_read)
  );
  assign io_halt = cpu_io_halt; // @[src/main/scala/cpu8086/CPU8086.scala 512:11]
  assign io_ax = cpu_io_ax; // @[src/main/scala/cpu8086/CPU8086.scala 513:9]
  assign io_bx = cpu_io_bx; // @[src/main/scala/cpu8086/CPU8086.scala 514:9]
  assign io_cx = cpu_io_cx; // @[src/main/scala/cpu8086/CPU8086.scala 515:9]
  assign io_dx = cpu_io_dx; // @[src/main/scala/cpu8086/CPU8086.scala 516:9]
  assign io_sp = cpu_io_sp; // @[src/main/scala/cpu8086/CPU8086.scala 517:9]
  assign io_ip = cpu_io_ip; // @[src/main/scala/cpu8086/CPU8086.scala 518:9]
  assign io_flags = cpu_io_flags; // @[src/main/scala/cpu8086/CPU8086.scala 519:12]
  assign cpu_clock = clock;
  assign cpu_reset = reset;
  assign cpu_io_memDataIn = mem_io_dataOut; // @[src/main/scala/cpu8086/CPU8086.scala 508:20]
  assign mem_clock = clock;
  assign mem_io_addr = cpu_io_memAddr; // @[src/main/scala/cpu8086/CPU8086.scala 506:15]
  assign mem_io_dataIn = cpu_io_memDataOut; // @[src/main/scala/cpu8086/CPU8086.scala 507:17]
  assign mem_io_write = cpu_io_memWrite; // @[src/main/scala/cpu8086/CPU8086.scala 509:16]
  assign mem_io_read = cpu_io_memRead; // @[src/main/scala/cpu8086/CPU8086.scala 510:15]
endmodule
